/*******************/
/* rom8x1024_sim.v */
/*******************/

//                  +----+
//  rom_addr[11:0]->|    |->rom_data[31:0]
//                  +----+

//
// ROM�ε��ҡ��������ߥ�졼������ѡ�
//

module rom8x1024_sim (rom_addr, rom_data);

  input   [11:0]  rom_addr;  // 12-bit ���ɥ쥹���ϥݡ���
  output  [31:0]  rom_data;  // 32-bit �ǡ������ϥݡ���

  reg     [31:0]  data;

  // Wire
  wire     [9:0]  word_addr; // 10-bit address, word

  assign word_addr = rom_addr[9:2];
   
  always @(word_addr) begin
    case (word_addr)
      10'h000: data = 32'he000001c; // 00400000: other type! opcode=56(10)
      10'h001: data = 32'h00000000; // 00400004: SLL, REG[0]<=REG[0]<<0;
      10'h002: data = 32'h00000000; // 00400008: SLL, REG[0]<=REG[0]<<0;
      10'h003: data = 32'h00000000; // 0040000c: SLL, REG[0]<=REG[0]<<0;
      10'h004: data = 32'h00000000; // 00400010: SLL, REG[0]<=REG[0]<<0;
      10'h005: data = 32'h00408950; // 00400014: R type, unknown. func=16(10)
      10'h006: data = 32'h00000000; // 00400018: SLL, REG[0]<=REG[0]<<0;
      10'h007: data = 32'h00000000; // 0040001c: SLL, REG[0]<=REG[0]<<0;
      10'h008: data = 32'h27bdffa8; // 00400020: ADDIU, REG[29]<=REG[29]+65448(=0x0000ffa8);
      10'h009: data = 32'hafbf0054; // 00400024: SW, RAM[REG[29]+84]<=REG[31];
      10'h00a: data = 32'hafbe0050; // 00400028: SW, RAM[REG[29]+80]<=REG[30];
      10'h00b: data = 32'h03a0f021; // 0040002c: ADDU, REG[30]<=REG[29]+REG[0];
      10'h00c: data = 32'h24020048; // 00400030: ADDIU, REG[2]<=REG[0]+72(=0x00000048);
      10'h00d: data = 32'hafc20010; // 00400034: SW, RAM[REG[30]+16]<=REG[2];
      10'h00e: data = 32'h24020045; // 00400038: ADDIU, REG[2]<=REG[0]+69(=0x00000045);
      10'h00f: data = 32'hafc20014; // 0040003c: SW, RAM[REG[30]+20]<=REG[2];
      10'h010: data = 32'h2402004c; // 00400040: ADDIU, REG[2]<=REG[0]+76(=0x0000004c);
      10'h011: data = 32'hafc20018; // 00400044: SW, RAM[REG[30]+24]<=REG[2];
      10'h012: data = 32'h2402004c; // 00400048: ADDIU, REG[2]<=REG[0]+76(=0x0000004c);
      10'h013: data = 32'hafc2001c; // 0040004c: SW, RAM[REG[30]+28]<=REG[2];
      10'h014: data = 32'h2402004f; // 00400050: ADDIU, REG[2]<=REG[0]+79(=0x0000004f);
      10'h015: data = 32'hafc20020; // 00400054: SW, RAM[REG[30]+32]<=REG[2];
      10'h016: data = 32'h2402000a; // 00400058: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h017: data = 32'hafc20024; // 0040005c: SW, RAM[REG[30]+36]<=REG[2];
      10'h018: data = 32'hafc00028; // 00400060: SW, RAM[REG[30]+40]<=REG[0];
      10'h019: data = 32'h27c20010; // 00400064: ADDIU, REG[2]<=REG[30]+16(=0x00000010);
      10'h01a: data = 32'h00402021; // 00400068: ADDU, REG[4]<=REG[2]+REG[0];
      10'h01b: data = 32'h0c10017e; // 0040006c: JAL, PC<=0x0010017e*4(=0x004005f8); REG[31]<=PC+4
      10'h01c: data = 32'h00000000; // 00400070: SLL, REG[0]<=REG[0]<<0;
      10'h01d: data = 32'h24020053; // 00400074: ADDIU, REG[2]<=REG[0]+83(=0x00000053);
      10'h01e: data = 32'hafc20010; // 00400078: SW, RAM[REG[30]+16]<=REG[2];
      10'h01f: data = 32'h24020054; // 0040007c: ADDIU, REG[2]<=REG[0]+84(=0x00000054);
      10'h020: data = 32'hafc20014; // 00400080: SW, RAM[REG[30]+20]<=REG[2];
      10'h021: data = 32'h24020052; // 00400084: ADDIU, REG[2]<=REG[0]+82(=0x00000052);
      10'h022: data = 32'hafc20018; // 00400088: SW, RAM[REG[30]+24]<=REG[2];
      10'h023: data = 32'h2402003d; // 0040008c: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h024: data = 32'hafc2001c; // 00400090: SW, RAM[REG[30]+28]<=REG[2];
      10'h025: data = 32'hafc00020; // 00400094: SW, RAM[REG[30]+32]<=REG[0];
      10'h026: data = 32'h27c20010; // 00400098: ADDIU, REG[2]<=REG[30]+16(=0x00000010);
      10'h027: data = 32'h00402021; // 0040009c: ADDU, REG[4]<=REG[2]+REG[0];
      10'h028: data = 32'h0c10017e; // 004000a0: JAL, PC<=0x0010017e*4(=0x004005f8); REG[31]<=PC+4
      10'h029: data = 32'h00000000; // 004000a4: SLL, REG[0]<=REG[0]<<0;
      10'h02a: data = 32'h0c10002e; // 004000a8: JAL, PC<=0x0010002e*4(=0x004000b8); REG[31]<=PC+4
      10'h02b: data = 32'h00000000; // 004000ac: SLL, REG[0]<=REG[0]<<0;
      10'h02c: data = 32'h0810001d; // 004000b0: J, PC<=0x0010001d*4(=0x00400074);
      10'h02d: data = 32'h00000000; // 004000b4: SLL, REG[0]<=REG[0]<<0;
      10'h02e: data = 32'h27bdff60; // 004000b8: ADDIU, REG[29]<=REG[29]+65376(=0x0000ff60);
      10'h02f: data = 32'hafbf009c; // 004000bc: SW, RAM[REG[29]+156]<=REG[31];
      10'h030: data = 32'hafbe0098; // 004000c0: SW, RAM[REG[29]+152]<=REG[30];
      10'h031: data = 32'h03a0f021; // 004000c4: ADDU, REG[30]<=REG[29]+REG[0];
      10'h032: data = 32'h27c20014; // 004000c8: ADDIU, REG[2]<=REG[30]+20(=0x00000014);
      10'h033: data = 32'h00402021; // 004000cc: ADDU, REG[4]<=REG[2]+REG[0];
      10'h034: data = 32'h0c10009c; // 004000d0: JAL, PC<=0x0010009c*4(=0x00400270); REG[31]<=PC+4
      10'h035: data = 32'h00000000; // 004000d4: SLL, REG[0]<=REG[0]<<0;
      10'h036: data = 32'hafc00010; // 004000d8: SW, RAM[REG[30]+16]<=REG[0];
      10'h037: data = 32'h08100049; // 004000dc: J, PC<=0x00100049*4(=0x00400124);
      10'h038: data = 32'h00000000; // 004000e0: SLL, REG[0]<=REG[0]<<0;
      10'h039: data = 32'h27c20014; // 004000e4: ADDIU, REG[2]<=REG[30]+20(=0x00000014);
      10'h03a: data = 32'h00402021; // 004000e8: ADDU, REG[4]<=REG[2]+REG[0];
      10'h03b: data = 32'h0c100061; // 004000ec: JAL, PC<=0x00100061*4(=0x00400184); REG[31]<=PC+4
      10'h03c: data = 32'h00000000; // 004000f0: SLL, REG[0]<=REG[0]<<0;
      10'h03d: data = 32'h10400005; // 004000f4: BEQ, PC<=(REG[2] == REG[0])?PC+4+5*4:PC+4;
      10'h03e: data = 32'h00000000; // 004000f8: SLL, REG[0]<=REG[0]<<0;
      10'h03f: data = 32'h0c100070; // 004000fc: JAL, PC<=0x00100070*4(=0x004001c0); REG[31]<=PC+4
      10'h040: data = 32'h00000000; // 00400100: SLL, REG[0]<=REG[0]<<0;
      10'h041: data = 32'h08100045; // 00400104: J, PC<=0x00100045*4(=0x00400114);
      10'h042: data = 32'h00000000; // 00400108: SLL, REG[0]<=REG[0]<<0;
      10'h043: data = 32'h0c100086; // 0040010c: JAL, PC<=0x00100086*4(=0x00400218); REG[31]<=PC+4
      10'h044: data = 32'h00000000; // 00400110: SLL, REG[0]<=REG[0]<<0;
      10'h045: data = 32'h8fc20010; // 00400114: LW, REG[2]<=RAM[REG[30]+16];
      10'h046: data = 32'h00000000; // 00400118: SLL, REG[0]<=REG[0]<<0;
      10'h047: data = 32'h24420001; // 0040011c: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h048: data = 32'hafc20010; // 00400120: SW, RAM[REG[30]+16]<=REG[2];
      10'h049: data = 32'h8fc20010; // 00400124: LW, REG[2]<=RAM[REG[30]+16];
      10'h04a: data = 32'h00000000; // 00400128: SLL, REG[0]<=REG[0]<<0;
      10'h04b: data = 32'h2c420101; // 0040012c: SLTIU, REG[2]<=(REG[2]<257(=0x00000101))?1:0;
      10'h04c: data = 32'h1440ffec; // 00400130: BNE, PC<=(REG[2] != REG[0])?PC+4+65516*4:PC+4;
      10'h04d: data = 32'h00000000; // 00400134: SLL, REG[0]<=REG[0]<<0;
      10'h04e: data = 32'h24020045; // 00400138: ADDIU, REG[2]<=REG[0]+69(=0x00000045);
      10'h04f: data = 32'hafc20054; // 0040013c: SW, RAM[REG[30]+84]<=REG[2];
      10'h050: data = 32'h2402004e; // 00400140: ADDIU, REG[2]<=REG[0]+78(=0x0000004e);
      10'h051: data = 32'hafc20058; // 00400144: SW, RAM[REG[30]+88]<=REG[2];
      10'h052: data = 32'h24020044; // 00400148: ADDIU, REG[2]<=REG[0]+68(=0x00000044);
      10'h053: data = 32'hafc2005c; // 0040014c: SW, RAM[REG[30]+92]<=REG[2];
      10'h054: data = 32'h2402000a; // 00400150: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h055: data = 32'hafc20060; // 00400154: SW, RAM[REG[30]+96]<=REG[2];
      10'h056: data = 32'hafc00064; // 00400158: SW, RAM[REG[30]+100]<=REG[0];
      10'h057: data = 32'h27c20054; // 0040015c: ADDIU, REG[2]<=REG[30]+84(=0x00000054);
      10'h058: data = 32'h00402021; // 00400160: ADDU, REG[4]<=REG[2]+REG[0];
      10'h059: data = 32'h0c10017e; // 00400164: JAL, PC<=0x0010017e*4(=0x004005f8); REG[31]<=PC+4
      10'h05a: data = 32'h00000000; // 00400168: SLL, REG[0]<=REG[0]<<0;
      10'h05b: data = 32'h03c0e821; // 0040016c: ADDU, REG[29]<=REG[30]+REG[0];
      10'h05c: data = 32'h8fbf009c; // 00400170: LW, REG[31]<=RAM[REG[29]+156];
      10'h05d: data = 32'h8fbe0098; // 00400174: LW, REG[30]<=RAM[REG[29]+152];
      10'h05e: data = 32'h27bd00a0; // 00400178: ADDIU, REG[29]<=REG[29]+160(=0x000000a0);
      10'h05f: data = 32'h03e00008; // 0040017c: JR, PC<=REG[31];
      10'h060: data = 32'h00000000; // 00400180: SLL, REG[0]<=REG[0]<<0;
      10'h061: data = 32'h27bdfff8; // 00400184: ADDIU, REG[29]<=REG[29]+65528(=0x0000fff8);
      10'h062: data = 32'hafbe0000; // 00400188: SW, RAM[REG[29]+0]<=REG[30];
      10'h063: data = 32'h03a0f021; // 0040018c: ADDU, REG[30]<=REG[29]+REG[0];
      10'h064: data = 32'hafc40008; // 00400190: SW, RAM[REG[30]+8]<=REG[4];
      10'h065: data = 32'h8fc20008; // 00400194: LW, REG[2]<=RAM[REG[30]+8];
      10'h066: data = 32'h00000000; // 00400198: SLL, REG[0]<=REG[0]<<0;
      10'h067: data = 32'h8c420000; // 0040019c: LW, REG[2]<=RAM[REG[2]+0];
      10'h068: data = 32'h00000000; // 004001a0: SLL, REG[0]<=REG[0]<<0;
      10'h069: data = 32'h3842004e; // 004001a4: XORI
      10'h06a: data = 32'h2c420001; // 004001a8: SLTIU, REG[2]<=(REG[2]<1(=0x00000001))?1:0;
      10'h06b: data = 32'h03c0e821; // 004001ac: ADDU, REG[29]<=REG[30]+REG[0];
      10'h06c: data = 32'h8fbe0000; // 004001b0: LW, REG[30]<=RAM[REG[29]+0];
      10'h06d: data = 32'h27bd0008; // 004001b4: ADDIU, REG[29]<=REG[29]+8(=0x00000008);
      10'h06e: data = 32'h03e00008; // 004001b8: JR, PC<=REG[31];
      10'h06f: data = 32'h00000000; // 004001bc: SLL, REG[0]<=REG[0]<<0;
      10'h070: data = 32'h27bdffe8; // 004001c0: ADDIU, REG[29]<=REG[29]+65512(=0x0000ffe8);
      10'h071: data = 32'hafbf0014; // 004001c4: SW, RAM[REG[29]+20]<=REG[31];
      10'h072: data = 32'hafbe0010; // 004001c8: SW, RAM[REG[29]+16]<=REG[30];
      10'h073: data = 32'h03a0f021; // 004001cc: ADDU, REG[30]<=REG[29]+REG[0];
      10'h074: data = 32'h24040008; // 004001d0: ADDIU, REG[4]<=REG[0]+8(=0x00000008);
      10'h075: data = 32'h0c10024b; // 004001d4: JAL, PC<=0x0010024b*4(=0x0040092c); REG[31]<=PC+4
      10'h076: data = 32'h00000000; // 004001d8: SLL, REG[0]<=REG[0]<<0;
      10'h077: data = 32'h24040004; // 004001dc: ADDIU, REG[4]<=REG[0]+4(=0x00000004);
      10'h078: data = 32'h0c10024b; // 004001e0: JAL, PC<=0x0010024b*4(=0x0040092c); REG[31]<=PC+4
      10'h079: data = 32'h00000000; // 004001e4: SLL, REG[0]<=REG[0]<<0;
      10'h07a: data = 32'h24040002; // 004001e8: ADDIU, REG[4]<=REG[0]+2(=0x00000002);
      10'h07b: data = 32'h0c10024b; // 004001ec: JAL, PC<=0x0010024b*4(=0x0040092c); REG[31]<=PC+4
      10'h07c: data = 32'h00000000; // 004001f0: SLL, REG[0]<=REG[0]<<0;
      10'h07d: data = 32'h24040001; // 004001f4: ADDIU, REG[4]<=REG[0]+1(=0x00000001);
      10'h07e: data = 32'h0c10024b; // 004001f8: JAL, PC<=0x0010024b*4(=0x0040092c); REG[31]<=PC+4
      10'h07f: data = 32'h00000000; // 004001fc: SLL, REG[0]<=REG[0]<<0;
      10'h080: data = 32'h03c0e821; // 00400200: ADDU, REG[29]<=REG[30]+REG[0];
      10'h081: data = 32'h8fbf0014; // 00400204: LW, REG[31]<=RAM[REG[29]+20];
      10'h082: data = 32'h8fbe0010; // 00400208: LW, REG[30]<=RAM[REG[29]+16];
      10'h083: data = 32'h27bd0018; // 0040020c: ADDIU, REG[29]<=REG[29]+24(=0x00000018);
      10'h084: data = 32'h03e00008; // 00400210: JR, PC<=REG[31];
      10'h085: data = 32'h00000000; // 00400214: SLL, REG[0]<=REG[0]<<0;
      10'h086: data = 32'h27bdffe8; // 00400218: ADDIU, REG[29]<=REG[29]+65512(=0x0000ffe8);
      10'h087: data = 32'hafbf0014; // 0040021c: SW, RAM[REG[29]+20]<=REG[31];
      10'h088: data = 32'hafbe0010; // 00400220: SW, RAM[REG[29]+16]<=REG[30];
      10'h089: data = 32'h03a0f021; // 00400224: ADDU, REG[30]<=REG[29]+REG[0];
      10'h08a: data = 32'h24040001; // 00400228: ADDIU, REG[4]<=REG[0]+1(=0x00000001);
      10'h08b: data = 32'h0c10024b; // 0040022c: JAL, PC<=0x0010024b*4(=0x0040092c); REG[31]<=PC+4
      10'h08c: data = 32'h00000000; // 00400230: SLL, REG[0]<=REG[0]<<0;
      10'h08d: data = 32'h24040002; // 00400234: ADDIU, REG[4]<=REG[0]+2(=0x00000002);
      10'h08e: data = 32'h0c10024b; // 00400238: JAL, PC<=0x0010024b*4(=0x0040092c); REG[31]<=PC+4
      10'h08f: data = 32'h00000000; // 0040023c: SLL, REG[0]<=REG[0]<<0;
      10'h090: data = 32'h24040004; // 00400240: ADDIU, REG[4]<=REG[0]+4(=0x00000004);
      10'h091: data = 32'h0c10024b; // 00400244: JAL, PC<=0x0010024b*4(=0x0040092c); REG[31]<=PC+4
      10'h092: data = 32'h00000000; // 00400248: SLL, REG[0]<=REG[0]<<0;
      10'h093: data = 32'h24040008; // 0040024c: ADDIU, REG[4]<=REG[0]+8(=0x00000008);
      10'h094: data = 32'h0c10024b; // 00400250: JAL, PC<=0x0010024b*4(=0x0040092c); REG[31]<=PC+4
      10'h095: data = 32'h00000000; // 00400254: SLL, REG[0]<=REG[0]<<0;
      10'h096: data = 32'h03c0e821; // 00400258: ADDU, REG[29]<=REG[30]+REG[0];
      10'h097: data = 32'h8fbf0014; // 0040025c: LW, REG[31]<=RAM[REG[29]+20];
      10'h098: data = 32'h8fbe0010; // 00400260: LW, REG[30]<=RAM[REG[29]+16];
      10'h099: data = 32'h27bd0018; // 00400264: ADDIU, REG[29]<=REG[29]+24(=0x00000018);
      10'h09a: data = 32'h03e00008; // 00400268: JR, PC<=REG[31];
      10'h09b: data = 32'h00000000; // 0040026c: SLL, REG[0]<=REG[0]<<0;
      10'h09c: data = 32'h27bdfff8; // 00400270: ADDIU, REG[29]<=REG[29]+65528(=0x0000fff8);
      10'h09d: data = 32'hafbe0000; // 00400274: SW, RAM[REG[29]+0]<=REG[30];
      10'h09e: data = 32'h03a0f021; // 00400278: ADDU, REG[30]<=REG[29]+REG[0];
      10'h09f: data = 32'hafc40008; // 0040027c: SW, RAM[REG[30]+8]<=REG[4];
      10'h0a0: data = 32'h24020308; // 00400280: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h0a1: data = 32'hac400000; // 00400284: SW, RAM[REG[2]+0]<=REG[0];
      10'h0a2: data = 32'h2403030c; // 00400288: ADDIU, REG[3]<=REG[0]+780(=0x0000030c);
      10'h0a3: data = 32'h24020001; // 0040028c: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h0a4: data = 32'hac620000; // 00400290: SW, RAM[REG[3]+0]<=REG[2];
      10'h0a5: data = 32'h24030308; // 00400294: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h0a6: data = 32'h24020001; // 00400298: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h0a7: data = 32'hac620000; // 0040029c: SW, RAM[REG[3]+0]<=REG[2];
      10'h0a8: data = 32'h24020308; // 004002a0: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h0a9: data = 32'hac400000; // 004002a4: SW, RAM[REG[2]+0]<=REG[0];
      10'h0aa: data = 32'h24030308; // 004002a8: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h0ab: data = 32'h24020001; // 004002ac: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h0ac: data = 32'hac620000; // 004002b0: SW, RAM[REG[3]+0]<=REG[2];
      10'h0ad: data = 32'h081000b4; // 004002b4: J, PC<=0x001000b4*4(=0x004002d0);
      10'h0ae: data = 32'h00000000; // 004002b8: SLL, REG[0]<=REG[0]<<0;
      10'h0af: data = 32'h24020308; // 004002bc: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h0b0: data = 32'hac400000; // 004002c0: SW, RAM[REG[2]+0]<=REG[0];
      10'h0b1: data = 32'h24030308; // 004002c4: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h0b2: data = 32'h24020001; // 004002c8: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h0b3: data = 32'hac620000; // 004002cc: SW, RAM[REG[3]+0]<=REG[2];
      10'h0b4: data = 32'h24020310; // 004002d0: ADDIU, REG[2]<=REG[0]+784(=0x00000310);
      10'h0b5: data = 32'h8c430000; // 004002d4: LW, REG[3]<=RAM[REG[2]+0];
      10'h0b6: data = 32'h2402ffff; // 004002d8: ADDIU, REG[2]<=REG[0]+65535(=0x0000ffff);
      10'h0b7: data = 32'h1062fff7; // 004002dc: BEQ, PC<=(REG[3] == REG[2])?PC+4+65527*4:PC+4;
      10'h0b8: data = 32'h00000000; // 004002e0: SLL, REG[0]<=REG[0]<<0;
      10'h0b9: data = 32'h08100162; // 004002e4: J, PC<=0x00100162*4(=0x00400588);
      10'h0ba: data = 32'h00000000; // 004002e8: SLL, REG[0]<=REG[0]<<0;
      10'h0bb: data = 32'h8fc20008; // 004002ec: LW, REG[2]<=RAM[REG[30]+8];
      10'h0bc: data = 32'h00000000; // 004002f0: SLL, REG[0]<=REG[0]<<0;
      10'h0bd: data = 32'h8c420000; // 004002f4: LW, REG[2]<=RAM[REG[2]+0];
      10'h0be: data = 32'h00000000; // 004002f8: SLL, REG[0]<=REG[0]<<0;
      10'h0bf: data = 32'h10400012; // 004002fc: BEQ, PC<=(REG[2] == REG[0])?PC+4+18*4:PC+4;
      10'h0c0: data = 32'h00000000; // 00400300: SLL, REG[0]<=REG[0]<<0;
      10'h0c1: data = 32'h8fc20008; // 00400304: LW, REG[2]<=RAM[REG[30]+8];
      10'h0c2: data = 32'h00000000; // 00400308: SLL, REG[0]<=REG[0]<<0;
      10'h0c3: data = 32'h8c420000; // 0040030c: LW, REG[2]<=RAM[REG[2]+0];
      10'h0c4: data = 32'h00000000; // 00400310: SLL, REG[0]<=REG[0]<<0;
      10'h0c5: data = 32'h2c42001b; // 00400314: SLTIU, REG[2]<=(REG[2]<27(=0x0000001b))?1:0;
      10'h0c6: data = 32'h1040000b; // 00400318: BEQ, PC<=(REG[2] == REG[0])?PC+4+11*4:PC+4;
      10'h0c7: data = 32'h00000000; // 0040031c: SLL, REG[0]<=REG[0]<<0;
      10'h0c8: data = 32'h8fc20008; // 00400320: LW, REG[2]<=RAM[REG[30]+8];
      10'h0c9: data = 32'h00000000; // 00400324: SLL, REG[0]<=REG[0]<<0;
      10'h0ca: data = 32'h8c420000; // 00400328: LW, REG[2]<=RAM[REG[2]+0];
      10'h0cb: data = 32'h00000000; // 0040032c: SLL, REG[0]<=REG[0]<<0;
      10'h0cc: data = 32'h24430040; // 00400330: ADDIU, REG[3]<=REG[2]+64(=0x00000040);
      10'h0cd: data = 32'h8fc20008; // 00400334: LW, REG[2]<=RAM[REG[30]+8];
      10'h0ce: data = 32'h00000000; // 00400338: SLL, REG[0]<=REG[0]<<0;
      10'h0cf: data = 32'hac430000; // 0040033c: SW, RAM[REG[2]+0]<=REG[3];
      10'h0d0: data = 32'h08100159; // 00400340: J, PC<=0x00100159*4(=0x00400564);
      10'h0d1: data = 32'h00000000; // 00400344: SLL, REG[0]<=REG[0]<<0;
      10'h0d2: data = 32'h8fc20008; // 00400348: LW, REG[2]<=RAM[REG[30]+8];
      10'h0d3: data = 32'h00000000; // 0040034c: SLL, REG[0]<=REG[0]<<0;
      10'h0d4: data = 32'h8c420000; // 00400350: LW, REG[2]<=RAM[REG[2]+0];
      10'h0d5: data = 32'h00000000; // 00400354: SLL, REG[0]<=REG[0]<<0;
      10'h0d6: data = 32'h2c420030; // 00400358: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h0d7: data = 32'h14400010; // 0040035c: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h0d8: data = 32'h00000000; // 00400360: SLL, REG[0]<=REG[0]<<0;
      10'h0d9: data = 32'h8fc20008; // 00400364: LW, REG[2]<=RAM[REG[30]+8];
      10'h0da: data = 32'h00000000; // 00400368: SLL, REG[0]<=REG[0]<<0;
      10'h0db: data = 32'h8c420000; // 0040036c: LW, REG[2]<=RAM[REG[2]+0];
      10'h0dc: data = 32'h00000000; // 00400370: SLL, REG[0]<=REG[0]<<0;
      10'h0dd: data = 32'h2c42003a; // 00400374: SLTIU, REG[2]<=(REG[2]<58(=0x0000003a))?1:0;
      10'h0de: data = 32'h10400009; // 00400378: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h0df: data = 32'h00000000; // 0040037c: SLL, REG[0]<=REG[0]<<0;
      10'h0e0: data = 32'h8fc20008; // 00400380: LW, REG[2]<=RAM[REG[30]+8];
      10'h0e1: data = 32'h00000000; // 00400384: SLL, REG[0]<=REG[0]<<0;
      10'h0e2: data = 32'h8c430000; // 00400388: LW, REG[3]<=RAM[REG[2]+0];
      10'h0e3: data = 32'h8fc20008; // 0040038c: LW, REG[2]<=RAM[REG[30]+8];
      10'h0e4: data = 32'h00000000; // 00400390: SLL, REG[0]<=REG[0]<<0;
      10'h0e5: data = 32'hac430000; // 00400394: SW, RAM[REG[2]+0]<=REG[3];
      10'h0e6: data = 32'h08100159; // 00400398: J, PC<=0x00100159*4(=0x00400564);
      10'h0e7: data = 32'h00000000; // 0040039c: SLL, REG[0]<=REG[0]<<0;
      10'h0e8: data = 32'h8fc20008; // 004003a0: LW, REG[2]<=RAM[REG[30]+8];
      10'h0e9: data = 32'h00000000; // 004003a4: SLL, REG[0]<=REG[0]<<0;
      10'h0ea: data = 32'h8c420000; // 004003a8: LW, REG[2]<=RAM[REG[2]+0];
      10'h0eb: data = 32'h00000000; // 004003ac: SLL, REG[0]<=REG[0]<<0;
      10'h0ec: data = 32'h14400006; // 004003b0: BNE, PC<=(REG[2] != REG[0])?PC+4+6*4:PC+4;
      10'h0ed: data = 32'h00000000; // 004003b4: SLL, REG[0]<=REG[0]<<0;
      10'h0ee: data = 32'h8fc30008; // 004003b8: LW, REG[3]<=RAM[REG[30]+8];
      10'h0ef: data = 32'h24020040; // 004003bc: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h0f0: data = 32'hac620000; // 004003c0: SW, RAM[REG[3]+0]<=REG[2];
      10'h0f1: data = 32'h08100159; // 004003c4: J, PC<=0x00100159*4(=0x00400564);
      10'h0f2: data = 32'h00000000; // 004003c8: SLL, REG[0]<=REG[0]<<0;
      10'h0f3: data = 32'h8fc20008; // 004003cc: LW, REG[2]<=RAM[REG[30]+8];
      10'h0f4: data = 32'h00000000; // 004003d0: SLL, REG[0]<=REG[0]<<0;
      10'h0f5: data = 32'h8c430000; // 004003d4: LW, REG[3]<=RAM[REG[2]+0];
      10'h0f6: data = 32'h2402001b; // 004003d8: ADDIU, REG[2]<=REG[0]+27(=0x0000001b);
      10'h0f7: data = 32'h14620006; // 004003dc: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0f8: data = 32'h00000000; // 004003e0: SLL, REG[0]<=REG[0]<<0;
      10'h0f9: data = 32'h8fc30008; // 004003e4: LW, REG[3]<=RAM[REG[30]+8];
      10'h0fa: data = 32'h2402005b; // 004003e8: ADDIU, REG[2]<=REG[0]+91(=0x0000005b);
      10'h0fb: data = 32'hac620000; // 004003ec: SW, RAM[REG[3]+0]<=REG[2];
      10'h0fc: data = 32'h08100159; // 004003f0: J, PC<=0x00100159*4(=0x00400564);
      10'h0fd: data = 32'h00000000; // 004003f4: SLL, REG[0]<=REG[0]<<0;
      10'h0fe: data = 32'h8fc20008; // 004003f8: LW, REG[2]<=RAM[REG[30]+8];
      10'h0ff: data = 32'h00000000; // 004003fc: SLL, REG[0]<=REG[0]<<0;
      10'h100: data = 32'h8c430000; // 00400400: LW, REG[3]<=RAM[REG[2]+0];
      10'h101: data = 32'h2402001d; // 00400404: ADDIU, REG[2]<=REG[0]+29(=0x0000001d);
      10'h102: data = 32'h14620006; // 00400408: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h103: data = 32'h00000000; // 0040040c: SLL, REG[0]<=REG[0]<<0;
      10'h104: data = 32'h8fc30008; // 00400410: LW, REG[3]<=RAM[REG[30]+8];
      10'h105: data = 32'h2402005d; // 00400414: ADDIU, REG[2]<=REG[0]+93(=0x0000005d);
      10'h106: data = 32'hac620000; // 00400418: SW, RAM[REG[3]+0]<=REG[2];
      10'h107: data = 32'h08100159; // 0040041c: J, PC<=0x00100159*4(=0x00400564);
      10'h108: data = 32'h00000000; // 00400420: SLL, REG[0]<=REG[0]<<0;
      10'h109: data = 32'h8fc20008; // 00400424: LW, REG[2]<=RAM[REG[30]+8];
      10'h10a: data = 32'h00000000; // 00400428: SLL, REG[0]<=REG[0]<<0;
      10'h10b: data = 32'h8c420000; // 0040042c: LW, REG[2]<=RAM[REG[2]+0];
      10'h10c: data = 32'h00000000; // 00400430: SLL, REG[0]<=REG[0]<<0;
      10'h10d: data = 32'h2c420020; // 00400434: SLTIU, REG[2]<=(REG[2]<32(=0x00000020))?1:0;
      10'h10e: data = 32'h14400010; // 00400438: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h10f: data = 32'h00000000; // 0040043c: SLL, REG[0]<=REG[0]<<0;
      10'h110: data = 32'h8fc20008; // 00400440: LW, REG[2]<=RAM[REG[30]+8];
      10'h111: data = 32'h00000000; // 00400444: SLL, REG[0]<=REG[0]<<0;
      10'h112: data = 32'h8c420000; // 00400448: LW, REG[2]<=RAM[REG[2]+0];
      10'h113: data = 32'h00000000; // 0040044c: SLL, REG[0]<=REG[0]<<0;
      10'h114: data = 32'h2c420030; // 00400450: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h115: data = 32'h10400009; // 00400454: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h116: data = 32'h00000000; // 00400458: SLL, REG[0]<=REG[0]<<0;
      10'h117: data = 32'h8fc20008; // 0040045c: LW, REG[2]<=RAM[REG[30]+8];
      10'h118: data = 32'h00000000; // 00400460: SLL, REG[0]<=REG[0]<<0;
      10'h119: data = 32'h8c430000; // 00400464: LW, REG[3]<=RAM[REG[2]+0];
      10'h11a: data = 32'h8fc20008; // 00400468: LW, REG[2]<=RAM[REG[30]+8];
      10'h11b: data = 32'h00000000; // 0040046c: SLL, REG[0]<=REG[0]<<0;
      10'h11c: data = 32'hac430000; // 00400470: SW, RAM[REG[2]+0]<=REG[3];
      10'h11d: data = 32'h08100159; // 00400474: J, PC<=0x00100159*4(=0x00400564);
      10'h11e: data = 32'h00000000; // 00400478: SLL, REG[0]<=REG[0]<<0;
      10'h11f: data = 32'h8fc20008; // 0040047c: LW, REG[2]<=RAM[REG[30]+8];
      10'h120: data = 32'h00000000; // 00400480: SLL, REG[0]<=REG[0]<<0;
      10'h121: data = 32'h8c430000; // 00400484: LW, REG[3]<=RAM[REG[2]+0];
      10'h122: data = 32'h2402003a; // 00400488: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h123: data = 32'h14620006; // 0040048c: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h124: data = 32'h00000000; // 00400490: SLL, REG[0]<=REG[0]<<0;
      10'h125: data = 32'h8fc30008; // 00400494: LW, REG[3]<=RAM[REG[30]+8];
      10'h126: data = 32'h2402003f; // 00400498: ADDIU, REG[2]<=REG[0]+63(=0x0000003f);
      10'h127: data = 32'hac620000; // 0040049c: SW, RAM[REG[3]+0]<=REG[2];
      10'h128: data = 32'h08100159; // 004004a0: J, PC<=0x00100159*4(=0x00400564);
      10'h129: data = 32'h00000000; // 004004a4: SLL, REG[0]<=REG[0]<<0;
      10'h12a: data = 32'h8fc20008; // 004004a8: LW, REG[2]<=RAM[REG[30]+8];
      10'h12b: data = 32'h00000000; // 004004ac: SLL, REG[0]<=REG[0]<<0;
      10'h12c: data = 32'h8c430000; // 004004b0: LW, REG[3]<=RAM[REG[2]+0];
      10'h12d: data = 32'h2402003b; // 004004b4: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h12e: data = 32'h14620006; // 004004b8: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h12f: data = 32'h00000000; // 004004bc: SLL, REG[0]<=REG[0]<<0;
      10'h130: data = 32'h8fc30008; // 004004c0: LW, REG[3]<=RAM[REG[30]+8];
      10'h131: data = 32'h2402003d; // 004004c4: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h132: data = 32'hac620000; // 004004c8: SW, RAM[REG[3]+0]<=REG[2];
      10'h133: data = 32'h08100159; // 004004cc: J, PC<=0x00100159*4(=0x00400564);
      10'h134: data = 32'h00000000; // 004004d0: SLL, REG[0]<=REG[0]<<0;
      10'h135: data = 32'h8fc20008; // 004004d4: LW, REG[2]<=RAM[REG[30]+8];
      10'h136: data = 32'h00000000; // 004004d8: SLL, REG[0]<=REG[0]<<0;
      10'h137: data = 32'h8c430000; // 004004dc: LW, REG[3]<=RAM[REG[2]+0];
      10'h138: data = 32'h2402003c; // 004004e0: ADDIU, REG[2]<=REG[0]+60(=0x0000003c);
      10'h139: data = 32'h14620006; // 004004e4: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h13a: data = 32'h00000000; // 004004e8: SLL, REG[0]<=REG[0]<<0;
      10'h13b: data = 32'h8fc30008; // 004004ec: LW, REG[3]<=RAM[REG[30]+8];
      10'h13c: data = 32'h2402003b; // 004004f0: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h13d: data = 32'hac620000; // 004004f4: SW, RAM[REG[3]+0]<=REG[2];
      10'h13e: data = 32'h08100159; // 004004f8: J, PC<=0x00100159*4(=0x00400564);
      10'h13f: data = 32'h00000000; // 004004fc: SLL, REG[0]<=REG[0]<<0;
      10'h140: data = 32'h8fc20008; // 00400500: LW, REG[2]<=RAM[REG[30]+8];
      10'h141: data = 32'h00000000; // 00400504: SLL, REG[0]<=REG[0]<<0;
      10'h142: data = 32'h8c430000; // 00400508: LW, REG[3]<=RAM[REG[2]+0];
      10'h143: data = 32'h2402003d; // 0040050c: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h144: data = 32'h14620006; // 00400510: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h145: data = 32'h00000000; // 00400514: SLL, REG[0]<=REG[0]<<0;
      10'h146: data = 32'h8fc30008; // 00400518: LW, REG[3]<=RAM[REG[30]+8];
      10'h147: data = 32'h2402003a; // 0040051c: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h148: data = 32'hac620000; // 00400520: SW, RAM[REG[3]+0]<=REG[2];
      10'h149: data = 32'h08100159; // 00400524: J, PC<=0x00100159*4(=0x00400564);
      10'h14a: data = 32'h00000000; // 00400528: SLL, REG[0]<=REG[0]<<0;
      10'h14b: data = 32'h8fc20008; // 0040052c: LW, REG[2]<=RAM[REG[30]+8];
      10'h14c: data = 32'h00000000; // 00400530: SLL, REG[0]<=REG[0]<<0;
      10'h14d: data = 32'h8c430000; // 00400534: LW, REG[3]<=RAM[REG[2]+0];
      10'h14e: data = 32'h2402003e; // 00400538: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h14f: data = 32'h14620006; // 0040053c: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h150: data = 32'h00000000; // 00400540: SLL, REG[0]<=REG[0]<<0;
      10'h151: data = 32'h8fc30008; // 00400544: LW, REG[3]<=RAM[REG[30]+8];
      10'h152: data = 32'h2402000a; // 00400548: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h153: data = 32'hac620000; // 0040054c: SW, RAM[REG[3]+0]<=REG[2];
      10'h154: data = 32'h08100159; // 00400550: J, PC<=0x00100159*4(=0x00400564);
      10'h155: data = 32'h00000000; // 00400554: SLL, REG[0]<=REG[0]<<0;
      10'h156: data = 32'h8fc30008; // 00400558: LW, REG[3]<=RAM[REG[30]+8];
      10'h157: data = 32'h24020040; // 0040055c: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h158: data = 32'hac620000; // 00400560: SW, RAM[REG[3]+0]<=REG[2];
      10'h159: data = 32'h24020308; // 00400564: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h15a: data = 32'hac400000; // 00400568: SW, RAM[REG[2]+0]<=REG[0];
      10'h15b: data = 32'h24030308; // 0040056c: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h15c: data = 32'h24020001; // 00400570: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h15d: data = 32'hac620000; // 00400574: SW, RAM[REG[3]+0]<=REG[2];
      10'h15e: data = 32'h8fc20008; // 00400578: LW, REG[2]<=RAM[REG[30]+8];
      10'h15f: data = 32'h00000000; // 0040057c: SLL, REG[0]<=REG[0]<<0;
      10'h160: data = 32'h24420004; // 00400580: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h161: data = 32'hafc20008; // 00400584: SW, RAM[REG[30]+8]<=REG[2];
      10'h162: data = 32'h24020310; // 00400588: ADDIU, REG[2]<=REG[0]+784(=0x00000310);
      10'h163: data = 32'h8c430000; // 0040058c: LW, REG[3]<=RAM[REG[2]+0];
      10'h164: data = 32'h8fc20008; // 00400590: LW, REG[2]<=RAM[REG[30]+8];
      10'h165: data = 32'h00000000; // 00400594: SLL, REG[0]<=REG[0]<<0;
      10'h166: data = 32'hac430000; // 00400598: SW, RAM[REG[2]+0]<=REG[3];
      10'h167: data = 32'h8fc20008; // 0040059c: LW, REG[2]<=RAM[REG[30]+8];
      10'h168: data = 32'h00000000; // 004005a0: SLL, REG[0]<=REG[0]<<0;
      10'h169: data = 32'h8c430000; // 004005a4: LW, REG[3]<=RAM[REG[2]+0];
      10'h16a: data = 32'h2402003e; // 004005a8: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h16b: data = 32'h1462ff4f; // 004005ac: BNE, PC<=(REG[3] != REG[2])?PC+4+65359*4:PC+4;
      10'h16c: data = 32'h00000000; // 004005b0: SLL, REG[0]<=REG[0]<<0;
      10'h16d: data = 32'h8fc20008; // 004005b4: LW, REG[2]<=RAM[REG[30]+8];
      10'h16e: data = 32'h00000000; // 004005b8: SLL, REG[0]<=REG[0]<<0;
      10'h16f: data = 32'hac400000; // 004005bc: SW, RAM[REG[2]+0]<=REG[0];
      10'h170: data = 32'h24020308; // 004005c0: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h171: data = 32'hac400000; // 004005c4: SW, RAM[REG[2]+0]<=REG[0];
      10'h172: data = 32'h2402030c; // 004005c8: ADDIU, REG[2]<=REG[0]+780(=0x0000030c);
      10'h173: data = 32'hac400000; // 004005cc: SW, RAM[REG[2]+0]<=REG[0];
      10'h174: data = 32'h24030308; // 004005d0: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h175: data = 32'h24020001; // 004005d4: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h176: data = 32'hac620000; // 004005d8: SW, RAM[REG[3]+0]<=REG[2];
      10'h177: data = 32'h24020308; // 004005dc: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h178: data = 32'hac400000; // 004005e0: SW, RAM[REG[2]+0]<=REG[0];
      10'h179: data = 32'h03c0e821; // 004005e4: ADDU, REG[29]<=REG[30]+REG[0];
      10'h17a: data = 32'h8fbe0000; // 004005e8: LW, REG[30]<=RAM[REG[29]+0];
      10'h17b: data = 32'h27bd0008; // 004005ec: ADDIU, REG[29]<=REG[29]+8(=0x00000008);
      10'h17c: data = 32'h03e00008; // 004005f0: JR, PC<=REG[31];
      10'h17d: data = 32'h00000000; // 004005f4: SLL, REG[0]<=REG[0]<<0;
      10'h17e: data = 32'h27bdfff8; // 004005f8: ADDIU, REG[29]<=REG[29]+65528(=0x0000fff8);
      10'h17f: data = 32'hafbe0000; // 004005fc: SW, RAM[REG[29]+0]<=REG[30];
      10'h180: data = 32'h03a0f021; // 00400600: ADDU, REG[30]<=REG[29]+REG[0];
      10'h181: data = 32'hafc40008; // 00400604: SW, RAM[REG[30]+8]<=REG[4];
      10'h182: data = 32'h08100240; // 00400608: J, PC<=0x00100240*4(=0x00400900);
      10'h183: data = 32'h00000000; // 0040060c: SLL, REG[0]<=REG[0]<<0;
      10'h184: data = 32'h24020300; // 00400610: ADDIU, REG[2]<=REG[0]+768(=0x00000300);
      10'h185: data = 32'hac400000; // 00400614: SW, RAM[REG[2]+0]<=REG[0];
      10'h186: data = 32'h8fc20008; // 00400618: LW, REG[2]<=RAM[REG[30]+8];
      10'h187: data = 32'h00000000; // 0040061c: SLL, REG[0]<=REG[0]<<0;
      10'h188: data = 32'h8c420000; // 00400620: LW, REG[2]<=RAM[REG[2]+0];
      10'h189: data = 32'h00000000; // 00400624: SLL, REG[0]<=REG[0]<<0;
      10'h18a: data = 32'h2c420041; // 00400628: SLTIU, REG[2]<=(REG[2]<65(=0x00000041))?1:0;
      10'h18b: data = 32'h14400011; // 0040062c: BNE, PC<=(REG[2] != REG[0])?PC+4+17*4:PC+4;
      10'h18c: data = 32'h00000000; // 00400630: SLL, REG[0]<=REG[0]<<0;
      10'h18d: data = 32'h8fc20008; // 00400634: LW, REG[2]<=RAM[REG[30]+8];
      10'h18e: data = 32'h00000000; // 00400638: SLL, REG[0]<=REG[0]<<0;
      10'h18f: data = 32'h8c420000; // 0040063c: LW, REG[2]<=RAM[REG[2]+0];
      10'h190: data = 32'h00000000; // 00400640: SLL, REG[0]<=REG[0]<<0;
      10'h191: data = 32'h2c42005b; // 00400644: SLTIU, REG[2]<=(REG[2]<91(=0x0000005b))?1:0;
      10'h192: data = 32'h1040000a; // 00400648: BEQ, PC<=(REG[2] == REG[0])?PC+4+10*4:PC+4;
      10'h193: data = 32'h00000000; // 0040064c: SLL, REG[0]<=REG[0]<<0;
      10'h194: data = 32'h24030304; // 00400650: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h195: data = 32'h8fc20008; // 00400654: LW, REG[2]<=RAM[REG[30]+8];
      10'h196: data = 32'h00000000; // 00400658: SLL, REG[0]<=REG[0]<<0;
      10'h197: data = 32'h8c420000; // 0040065c: LW, REG[2]<=RAM[REG[2]+0];
      10'h198: data = 32'h00000000; // 00400660: SLL, REG[0]<=REG[0]<<0;
      10'h199: data = 32'h2442ffc0; // 00400664: ADDIU, REG[2]<=REG[2]+65472(=0x0000ffc0);
      10'h19a: data = 32'hac620000; // 00400668: SW, RAM[REG[3]+0]<=REG[2];
      10'h19b: data = 32'h08100239; // 0040066c: J, PC<=0x00100239*4(=0x004008e4);
      10'h19c: data = 32'h00000000; // 00400670: SLL, REG[0]<=REG[0]<<0;
      10'h19d: data = 32'h8fc20008; // 00400674: LW, REG[2]<=RAM[REG[30]+8];
      10'h19e: data = 32'h00000000; // 00400678: SLL, REG[0]<=REG[0]<<0;
      10'h19f: data = 32'h8c420000; // 0040067c: LW, REG[2]<=RAM[REG[2]+0];
      10'h1a0: data = 32'h00000000; // 00400680: SLL, REG[0]<=REG[0]<<0;
      10'h1a1: data = 32'h2c420061; // 00400684: SLTIU, REG[2]<=(REG[2]<97(=0x00000061))?1:0;
      10'h1a2: data = 32'h14400011; // 00400688: BNE, PC<=(REG[2] != REG[0])?PC+4+17*4:PC+4;
      10'h1a3: data = 32'h00000000; // 0040068c: SLL, REG[0]<=REG[0]<<0;
      10'h1a4: data = 32'h8fc20008; // 00400690: LW, REG[2]<=RAM[REG[30]+8];
      10'h1a5: data = 32'h00000000; // 00400694: SLL, REG[0]<=REG[0]<<0;
      10'h1a6: data = 32'h8c420000; // 00400698: LW, REG[2]<=RAM[REG[2]+0];
      10'h1a7: data = 32'h00000000; // 0040069c: SLL, REG[0]<=REG[0]<<0;
      10'h1a8: data = 32'h2c42007b; // 004006a0: SLTIU, REG[2]<=(REG[2]<123(=0x0000007b))?1:0;
      10'h1a9: data = 32'h1040000a; // 004006a4: BEQ, PC<=(REG[2] == REG[0])?PC+4+10*4:PC+4;
      10'h1aa: data = 32'h00000000; // 004006a8: SLL, REG[0]<=REG[0]<<0;
      10'h1ab: data = 32'h24030304; // 004006ac: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h1ac: data = 32'h8fc20008; // 004006b0: LW, REG[2]<=RAM[REG[30]+8];
      10'h1ad: data = 32'h00000000; // 004006b4: SLL, REG[0]<=REG[0]<<0;
      10'h1ae: data = 32'h8c420000; // 004006b8: LW, REG[2]<=RAM[REG[2]+0];
      10'h1af: data = 32'h00000000; // 004006bc: SLL, REG[0]<=REG[0]<<0;
      10'h1b0: data = 32'h2442ffa0; // 004006c0: ADDIU, REG[2]<=REG[2]+65440(=0x0000ffa0);
      10'h1b1: data = 32'hac620000; // 004006c4: SW, RAM[REG[3]+0]<=REG[2];
      10'h1b2: data = 32'h08100239; // 004006c8: J, PC<=0x00100239*4(=0x004008e4);
      10'h1b3: data = 32'h00000000; // 004006cc: SLL, REG[0]<=REG[0]<<0;
      10'h1b4: data = 32'h8fc20008; // 004006d0: LW, REG[2]<=RAM[REG[30]+8];
      10'h1b5: data = 32'h00000000; // 004006d4: SLL, REG[0]<=REG[0]<<0;
      10'h1b6: data = 32'h8c420000; // 004006d8: LW, REG[2]<=RAM[REG[2]+0];
      10'h1b7: data = 32'h00000000; // 004006dc: SLL, REG[0]<=REG[0]<<0;
      10'h1b8: data = 32'h2c420030; // 004006e0: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h1b9: data = 32'h14400010; // 004006e4: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h1ba: data = 32'h00000000; // 004006e8: SLL, REG[0]<=REG[0]<<0;
      10'h1bb: data = 32'h8fc20008; // 004006ec: LW, REG[2]<=RAM[REG[30]+8];
      10'h1bc: data = 32'h00000000; // 004006f0: SLL, REG[0]<=REG[0]<<0;
      10'h1bd: data = 32'h8c420000; // 004006f4: LW, REG[2]<=RAM[REG[2]+0];
      10'h1be: data = 32'h00000000; // 004006f8: SLL, REG[0]<=REG[0]<<0;
      10'h1bf: data = 32'h2c42003a; // 004006fc: SLTIU, REG[2]<=(REG[2]<58(=0x0000003a))?1:0;
      10'h1c0: data = 32'h10400009; // 00400700: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h1c1: data = 32'h00000000; // 00400704: SLL, REG[0]<=REG[0]<<0;
      10'h1c2: data = 32'h24020304; // 00400708: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h1c3: data = 32'h8fc30008; // 0040070c: LW, REG[3]<=RAM[REG[30]+8];
      10'h1c4: data = 32'h00000000; // 00400710: SLL, REG[0]<=REG[0]<<0;
      10'h1c5: data = 32'h8c630000; // 00400714: LW, REG[3]<=RAM[REG[3]+0];
      10'h1c6: data = 32'h00000000; // 00400718: SLL, REG[0]<=REG[0]<<0;
      10'h1c7: data = 32'hac430000; // 0040071c: SW, RAM[REG[2]+0]<=REG[3];
      10'h1c8: data = 32'h08100239; // 00400720: J, PC<=0x00100239*4(=0x004008e4);
      10'h1c9: data = 32'h00000000; // 00400724: SLL, REG[0]<=REG[0]<<0;
      10'h1ca: data = 32'h8fc20008; // 00400728: LW, REG[2]<=RAM[REG[30]+8];
      10'h1cb: data = 32'h00000000; // 0040072c: SLL, REG[0]<=REG[0]<<0;
      10'h1cc: data = 32'h8c430000; // 00400730: LW, REG[3]<=RAM[REG[2]+0];
      10'h1cd: data = 32'h24020040; // 00400734: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h1ce: data = 32'h14620005; // 00400738: BNE, PC<=(REG[3] != REG[2])?PC+4+5*4:PC+4;
      10'h1cf: data = 32'h00000000; // 0040073c: SLL, REG[0]<=REG[0]<<0;
      10'h1d0: data = 32'h24020304; // 00400740: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h1d1: data = 32'hac400000; // 00400744: SW, RAM[REG[2]+0]<=REG[0];
      10'h1d2: data = 32'h08100239; // 00400748: J, PC<=0x00100239*4(=0x004008e4);
      10'h1d3: data = 32'h00000000; // 0040074c: SLL, REG[0]<=REG[0]<<0;
      10'h1d4: data = 32'h8fc20008; // 00400750: LW, REG[2]<=RAM[REG[30]+8];
      10'h1d5: data = 32'h00000000; // 00400754: SLL, REG[0]<=REG[0]<<0;
      10'h1d6: data = 32'h8c430000; // 00400758: LW, REG[3]<=RAM[REG[2]+0];
      10'h1d7: data = 32'h2402005b; // 0040075c: ADDIU, REG[2]<=REG[0]+91(=0x0000005b);
      10'h1d8: data = 32'h14620006; // 00400760: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h1d9: data = 32'h00000000; // 00400764: SLL, REG[0]<=REG[0]<<0;
      10'h1da: data = 32'h24030304; // 00400768: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h1db: data = 32'h2402001b; // 0040076c: ADDIU, REG[2]<=REG[0]+27(=0x0000001b);
      10'h1dc: data = 32'hac620000; // 00400770: SW, RAM[REG[3]+0]<=REG[2];
      10'h1dd: data = 32'h08100239; // 00400774: J, PC<=0x00100239*4(=0x004008e4);
      10'h1de: data = 32'h00000000; // 00400778: SLL, REG[0]<=REG[0]<<0;
      10'h1df: data = 32'h8fc20008; // 0040077c: LW, REG[2]<=RAM[REG[30]+8];
      10'h1e0: data = 32'h00000000; // 00400780: SLL, REG[0]<=REG[0]<<0;
      10'h1e1: data = 32'h8c430000; // 00400784: LW, REG[3]<=RAM[REG[2]+0];
      10'h1e2: data = 32'h2402005d; // 00400788: ADDIU, REG[2]<=REG[0]+93(=0x0000005d);
      10'h1e3: data = 32'h14620006; // 0040078c: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h1e4: data = 32'h00000000; // 00400790: SLL, REG[0]<=REG[0]<<0;
      10'h1e5: data = 32'h24030304; // 00400794: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h1e6: data = 32'h2402001d; // 00400798: ADDIU, REG[2]<=REG[0]+29(=0x0000001d);
      10'h1e7: data = 32'hac620000; // 0040079c: SW, RAM[REG[3]+0]<=REG[2];
      10'h1e8: data = 32'h08100239; // 004007a0: J, PC<=0x00100239*4(=0x004008e4);
      10'h1e9: data = 32'h00000000; // 004007a4: SLL, REG[0]<=REG[0]<<0;
      10'h1ea: data = 32'h8fc20008; // 004007a8: LW, REG[2]<=RAM[REG[30]+8];
      10'h1eb: data = 32'h00000000; // 004007ac: SLL, REG[0]<=REG[0]<<0;
      10'h1ec: data = 32'h8c420000; // 004007b0: LW, REG[2]<=RAM[REG[2]+0];
      10'h1ed: data = 32'h00000000; // 004007b4: SLL, REG[0]<=REG[0]<<0;
      10'h1ee: data = 32'h2c420020; // 004007b8: SLTIU, REG[2]<=(REG[2]<32(=0x00000020))?1:0;
      10'h1ef: data = 32'h14400010; // 004007bc: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h1f0: data = 32'h00000000; // 004007c0: SLL, REG[0]<=REG[0]<<0;
      10'h1f1: data = 32'h8fc20008; // 004007c4: LW, REG[2]<=RAM[REG[30]+8];
      10'h1f2: data = 32'h00000000; // 004007c8: SLL, REG[0]<=REG[0]<<0;
      10'h1f3: data = 32'h8c420000; // 004007cc: LW, REG[2]<=RAM[REG[2]+0];
      10'h1f4: data = 32'h00000000; // 004007d0: SLL, REG[0]<=REG[0]<<0;
      10'h1f5: data = 32'h2c420030; // 004007d4: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h1f6: data = 32'h10400009; // 004007d8: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h1f7: data = 32'h00000000; // 004007dc: SLL, REG[0]<=REG[0]<<0;
      10'h1f8: data = 32'h24020304; // 004007e0: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h1f9: data = 32'h8fc30008; // 004007e4: LW, REG[3]<=RAM[REG[30]+8];
      10'h1fa: data = 32'h00000000; // 004007e8: SLL, REG[0]<=REG[0]<<0;
      10'h1fb: data = 32'h8c630000; // 004007ec: LW, REG[3]<=RAM[REG[3]+0];
      10'h1fc: data = 32'h00000000; // 004007f0: SLL, REG[0]<=REG[0]<<0;
      10'h1fd: data = 32'hac430000; // 004007f4: SW, RAM[REG[2]+0]<=REG[3];
      10'h1fe: data = 32'h08100239; // 004007f8: J, PC<=0x00100239*4(=0x004008e4);
      10'h1ff: data = 32'h00000000; // 004007fc: SLL, REG[0]<=REG[0]<<0;
      10'h200: data = 32'h8fc20008; // 00400800: LW, REG[2]<=RAM[REG[30]+8];
      10'h201: data = 32'h00000000; // 00400804: SLL, REG[0]<=REG[0]<<0;
      10'h202: data = 32'h8c430000; // 00400808: LW, REG[3]<=RAM[REG[2]+0];
      10'h203: data = 32'h2402003f; // 0040080c: ADDIU, REG[2]<=REG[0]+63(=0x0000003f);
      10'h204: data = 32'h14620006; // 00400810: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h205: data = 32'h00000000; // 00400814: SLL, REG[0]<=REG[0]<<0;
      10'h206: data = 32'h24030304; // 00400818: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h207: data = 32'h2402003a; // 0040081c: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h208: data = 32'hac620000; // 00400820: SW, RAM[REG[3]+0]<=REG[2];
      10'h209: data = 32'h08100239; // 00400824: J, PC<=0x00100239*4(=0x004008e4);
      10'h20a: data = 32'h00000000; // 00400828: SLL, REG[0]<=REG[0]<<0;
      10'h20b: data = 32'h8fc20008; // 0040082c: LW, REG[2]<=RAM[REG[30]+8];
      10'h20c: data = 32'h00000000; // 00400830: SLL, REG[0]<=REG[0]<<0;
      10'h20d: data = 32'h8c430000; // 00400834: LW, REG[3]<=RAM[REG[2]+0];
      10'h20e: data = 32'h2402003d; // 00400838: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h20f: data = 32'h14620006; // 0040083c: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h210: data = 32'h00000000; // 00400840: SLL, REG[0]<=REG[0]<<0;
      10'h211: data = 32'h24030304; // 00400844: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h212: data = 32'h2402003b; // 00400848: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h213: data = 32'hac620000; // 0040084c: SW, RAM[REG[3]+0]<=REG[2];
      10'h214: data = 32'h08100239; // 00400850: J, PC<=0x00100239*4(=0x004008e4);
      10'h215: data = 32'h00000000; // 00400854: SLL, REG[0]<=REG[0]<<0;
      10'h216: data = 32'h8fc20008; // 00400858: LW, REG[2]<=RAM[REG[30]+8];
      10'h217: data = 32'h00000000; // 0040085c: SLL, REG[0]<=REG[0]<<0;
      10'h218: data = 32'h8c430000; // 00400860: LW, REG[3]<=RAM[REG[2]+0];
      10'h219: data = 32'h2402003b; // 00400864: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h21a: data = 32'h14620006; // 00400868: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h21b: data = 32'h00000000; // 0040086c: SLL, REG[0]<=REG[0]<<0;
      10'h21c: data = 32'h24030304; // 00400870: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h21d: data = 32'h2402003c; // 00400874: ADDIU, REG[2]<=REG[0]+60(=0x0000003c);
      10'h21e: data = 32'hac620000; // 00400878: SW, RAM[REG[3]+0]<=REG[2];
      10'h21f: data = 32'h08100239; // 0040087c: J, PC<=0x00100239*4(=0x004008e4);
      10'h220: data = 32'h00000000; // 00400880: SLL, REG[0]<=REG[0]<<0;
      10'h221: data = 32'h8fc20008; // 00400884: LW, REG[2]<=RAM[REG[30]+8];
      10'h222: data = 32'h00000000; // 00400888: SLL, REG[0]<=REG[0]<<0;
      10'h223: data = 32'h8c430000; // 0040088c: LW, REG[3]<=RAM[REG[2]+0];
      10'h224: data = 32'h2402003a; // 00400890: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h225: data = 32'h14620006; // 00400894: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h226: data = 32'h00000000; // 00400898: SLL, REG[0]<=REG[0]<<0;
      10'h227: data = 32'h24030304; // 0040089c: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h228: data = 32'h2402003d; // 004008a0: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h229: data = 32'hac620000; // 004008a4: SW, RAM[REG[3]+0]<=REG[2];
      10'h22a: data = 32'h08100239; // 004008a8: J, PC<=0x00100239*4(=0x004008e4);
      10'h22b: data = 32'h00000000; // 004008ac: SLL, REG[0]<=REG[0]<<0;
      10'h22c: data = 32'h8fc20008; // 004008b0: LW, REG[2]<=RAM[REG[30]+8];
      10'h22d: data = 32'h00000000; // 004008b4: SLL, REG[0]<=REG[0]<<0;
      10'h22e: data = 32'h8c430000; // 004008b8: LW, REG[3]<=RAM[REG[2]+0];
      10'h22f: data = 32'h2402000a; // 004008bc: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h230: data = 32'h14620006; // 004008c0: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h231: data = 32'h00000000; // 004008c4: SLL, REG[0]<=REG[0]<<0;
      10'h232: data = 32'h24030304; // 004008c8: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h233: data = 32'h2402003e; // 004008cc: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h234: data = 32'hac620000; // 004008d0: SW, RAM[REG[3]+0]<=REG[2];
      10'h235: data = 32'h08100239; // 004008d4: J, PC<=0x00100239*4(=0x004008e4);
      10'h236: data = 32'h00000000; // 004008d8: SLL, REG[0]<=REG[0]<<0;
      10'h237: data = 32'h24020304; // 004008dc: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h238: data = 32'hac400000; // 004008e0: SW, RAM[REG[2]+0]<=REG[0];
      10'h239: data = 32'h24030300; // 004008e4: ADDIU, REG[3]<=REG[0]+768(=0x00000300);
      10'h23a: data = 32'h24020001; // 004008e8: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h23b: data = 32'hac620000; // 004008ec: SW, RAM[REG[3]+0]<=REG[2];
      10'h23c: data = 32'h8fc20008; // 004008f0: LW, REG[2]<=RAM[REG[30]+8];
      10'h23d: data = 32'h00000000; // 004008f4: SLL, REG[0]<=REG[0]<<0;
      10'h23e: data = 32'h24420004; // 004008f8: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h23f: data = 32'hafc20008; // 004008fc: SW, RAM[REG[30]+8]<=REG[2];
      10'h240: data = 32'h8fc20008; // 00400900: LW, REG[2]<=RAM[REG[30]+8];
      10'h241: data = 32'h00000000; // 00400904: SLL, REG[0]<=REG[0]<<0;
      10'h242: data = 32'h8c420000; // 00400908: LW, REG[2]<=RAM[REG[2]+0];
      10'h243: data = 32'h00000000; // 0040090c: SLL, REG[0]<=REG[0]<<0;
      10'h244: data = 32'h1440ff3f; // 00400910: BNE, PC<=(REG[2] != REG[0])?PC+4+65343*4:PC+4;
      10'h245: data = 32'h00000000; // 00400914: SLL, REG[0]<=REG[0]<<0;
      10'h246: data = 32'h03c0e821; // 00400918: ADDU, REG[29]<=REG[30]+REG[0];
      10'h247: data = 32'h8fbe0000; // 0040091c: LW, REG[30]<=RAM[REG[29]+0];
      10'h248: data = 32'h27bd0008; // 00400920: ADDIU, REG[29]<=REG[29]+8(=0x00000008);
      10'h249: data = 32'h03e00008; // 00400924: JR, PC<=REG[31];
      10'h24a: data = 32'h00000000; // 00400928: SLL, REG[0]<=REG[0]<<0;
      10'h24b: data = 32'h27bdfff0; // 0040092c: ADDIU, REG[29]<=REG[29]+65520(=0x0000fff0);
      10'h24c: data = 32'hafbe0008; // 00400930: SW, RAM[REG[29]+8]<=REG[30];
      10'h24d: data = 32'h03a0f021; // 00400934: ADDU, REG[30]<=REG[29]+REG[0];
      10'h24e: data = 32'hafc40010; // 00400938: SW, RAM[REG[30]+16]<=REG[4];
      10'h24f: data = 32'h24030320; // 0040093c: ADDIU, REG[3]<=REG[0]+800(=0x00000320);
      10'h250: data = 32'h8fc20010; // 00400940: LW, REG[2]<=RAM[REG[30]+16];
      10'h251: data = 32'h00000000; // 00400944: SLL, REG[0]<=REG[0]<<0;
      10'h252: data = 32'hac620000; // 00400948: SW, RAM[REG[3]+0]<=REG[2];
      10'h253: data = 32'h03c0e821; // 0040094c: ADDU, REG[29]<=REG[30]+REG[0];
      10'h254: data = 32'h8fbe0008; // 00400950: LW, REG[30]<=RAM[REG[29]+8];
      10'h255: data = 32'h27bd0010; // 00400954: ADDIU, REG[29]<=REG[29]+16(=0x00000010);
      10'h256: data = 32'h03e00008; // 00400958: JR, PC<=REG[31];
      10'h257: data = 32'h00000000; // 0040095c: SLL, REG[0]<=REG[0]<<0;
    endcase
  end

  assign rom_data = data;
endmodule
