/*******************/
/* rom8x1024_sim.v */
/*******************/

//                  +----+
//  rom_addr[11:0]->|    |->rom_data[31:0]
//                  +----+

//
// ROM�ε��ҡ��������ߥ�졼������ѡ�
//

module rom8x1024_sim (rom_addr, rom_data);

  input   [11:0]  rom_addr;  // 12-bit ���ɥ쥹���ϥݡ���
  output  [31:0]  rom_data;  // 32-bit �ǡ������ϥݡ���

  reg     [31:0]  data;

  // Wire
  wire     [9:0]  word_addr; // 10-bit address, word

  assign word_addr = rom_addr[9:2];
   
  always @(word_addr) begin
    case (word_addr)
      10'h000: data = 32'he000001c; // 00400000: other type! opcode=56(10)
      10'h001: data = 32'h00000000; // 00400004: SLL, REG[0]<=REG[0]<<0;
      10'h002: data = 32'h00000000; // 00400008: SLL, REG[0]<=REG[0]<<0;
      10'h003: data = 32'h00000000; // 0040000c: SLL, REG[0]<=REG[0]<<0;
      10'h004: data = 32'h00000000; // 00400010: SLL, REG[0]<=REG[0]<<0;
      10'h005: data = 32'h00408930; // 00400014: R type, unknown. func=48(10)
      10'h006: data = 32'h00000000; // 00400018: SLL, REG[0]<=REG[0]<<0;
      10'h007: data = 32'h00000000; // 0040001c: SLL, REG[0]<=REG[0]<<0;
      10'h008: data = 32'h27bdffa8; // 00400020: ADDIU, REG[29]<=REG[29]+65448(=0x0000ffa8);
      10'h009: data = 32'hafbf0054; // 00400024: SW, RAM[REG[29]+84]<=REG[31];
      10'h00a: data = 32'hafbe0050; // 00400028: SW, RAM[REG[29]+80]<=REG[30];
      10'h00b: data = 32'h03a0f021; // 0040002c: ADDU, REG[30]<=REG[29]+REG[0];
      10'h00c: data = 32'h24020048; // 00400030: ADDIU, REG[2]<=REG[0]+72(=0x00000048);
      10'h00d: data = 32'hafc20010; // 00400034: SW, RAM[REG[30]+16]<=REG[2];
      10'h00e: data = 32'h24020045; // 00400038: ADDIU, REG[2]<=REG[0]+69(=0x00000045);
      10'h00f: data = 32'hafc20014; // 0040003c: SW, RAM[REG[30]+20]<=REG[2];
      10'h010: data = 32'h2402004c; // 00400040: ADDIU, REG[2]<=REG[0]+76(=0x0000004c);
      10'h011: data = 32'hafc20018; // 00400044: SW, RAM[REG[30]+24]<=REG[2];
      10'h012: data = 32'h2402004c; // 00400048: ADDIU, REG[2]<=REG[0]+76(=0x0000004c);
      10'h013: data = 32'hafc2001c; // 0040004c: SW, RAM[REG[30]+28]<=REG[2];
      10'h014: data = 32'h2402004f; // 00400050: ADDIU, REG[2]<=REG[0]+79(=0x0000004f);
      10'h015: data = 32'hafc20020; // 00400054: SW, RAM[REG[30]+32]<=REG[2];
      10'h016: data = 32'h2402000a; // 00400058: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h017: data = 32'hafc20024; // 0040005c: SW, RAM[REG[30]+36]<=REG[2];
      10'h018: data = 32'hafc00028; // 00400060: SW, RAM[REG[30]+40]<=REG[0];
      10'h019: data = 32'h27c20010; // 00400064: ADDIU, REG[2]<=REG[30]+16(=0x00000010);
      10'h01a: data = 32'h00402021; // 00400068: ADDU, REG[4]<=REG[2]+REG[0];
      10'h01b: data = 32'h0c100174; // 0040006c: JAL, PC<=0x00100174*4(=0x004005d0); REG[31]<=PC+4
      10'h01c: data = 32'h00000000; // 00400070: SLL, REG[0]<=REG[0]<<0;
      10'h01d: data = 32'h2402004e; // 00400074: ADDIU, REG[2]<=REG[0]+78(=0x0000004e);
      10'h01e: data = 32'hafc20010; // 00400078: SW, RAM[REG[30]+16]<=REG[2];
      10'h01f: data = 32'h24020055; // 0040007c: ADDIU, REG[2]<=REG[0]+85(=0x00000055);
      10'h020: data = 32'hafc20014; // 00400080: SW, RAM[REG[30]+20]<=REG[2];
      10'h021: data = 32'h2402004d; // 00400084: ADDIU, REG[2]<=REG[0]+77(=0x0000004d);
      10'h022: data = 32'hafc20018; // 00400088: SW, RAM[REG[30]+24]<=REG[2];
      10'h023: data = 32'h2402003d; // 0040008c: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h024: data = 32'hafc2001c; // 00400090: SW, RAM[REG[30]+28]<=REG[2];
      10'h025: data = 32'hafc00020; // 00400094: SW, RAM[REG[30]+32]<=REG[0];
      10'h026: data = 32'h27c20010; // 00400098: ADDIU, REG[2]<=REG[30]+16(=0x00000010);
      10'h027: data = 32'h00402021; // 0040009c: ADDU, REG[4]<=REG[2]+REG[0];
      10'h028: data = 32'h0c100174; // 004000a0: JAL, PC<=0x00100174*4(=0x004005d0); REG[31]<=PC+4
      10'h029: data = 32'h00000000; // 004000a4: SLL, REG[0]<=REG[0]<<0;
      10'h02a: data = 32'h0c10002e; // 004000a8: JAL, PC<=0x0010002e*4(=0x004000b8); REG[31]<=PC+4
      10'h02b: data = 32'h00000000; // 004000ac: SLL, REG[0]<=REG[0]<<0;
      10'h02c: data = 32'h0810001d; // 004000b0: J, PC<=0x0010001d*4(=0x00400074);
      10'h02d: data = 32'h00000000; // 004000b4: SLL, REG[0]<=REG[0]<<0;
      10'h02e: data = 32'h27bdffa0; // 004000b8: ADDIU, REG[29]<=REG[29]+65440(=0x0000ffa0);
      10'h02f: data = 32'hafbf005c; // 004000bc: SW, RAM[REG[29]+92]<=REG[31];
      10'h030: data = 32'hafbe0058; // 004000c0: SW, RAM[REG[29]+88]<=REG[30];
      10'h031: data = 32'h03a0f021; // 004000c4: ADDU, REG[30]<=REG[29]+REG[0];
      10'h032: data = 32'h27c20014; // 004000c8: ADDIU, REG[2]<=REG[30]+20(=0x00000014);
      10'h033: data = 32'h00402021; // 004000cc: ADDU, REG[4]<=REG[2]+REG[0];
      10'h034: data = 32'h0c100092; // 004000d0: JAL, PC<=0x00100092*4(=0x00400248); REG[31]<=PC+4
      10'h035: data = 32'h00000000; // 004000d4: SLL, REG[0]<=REG[0]<<0;
      10'h036: data = 32'hafc00010; // 004000d8: SW, RAM[REG[30]+16]<=REG[0];
      10'h037: data = 32'h0810004c; // 004000dc: J, PC<=0x0010004c*4(=0x00400130);
      10'h038: data = 32'h00000000; // 004000e0: SLL, REG[0]<=REG[0]<<0;
      10'h039: data = 32'h27c20014; // 004000e4: ADDIU, REG[2]<=REG[30]+20(=0x00000014);
      10'h03a: data = 32'h00402021; // 004000e8: ADDU, REG[4]<=REG[2]+REG[0];
      10'h03b: data = 32'h0c100057; // 004000ec: JAL, PC<=0x00100057*4(=0x0040015c); REG[31]<=PC+4
      10'h03c: data = 32'h00000000; // 004000f0: SLL, REG[0]<=REG[0]<<0;
      10'h03d: data = 32'h10400008; // 004000f4: BEQ, PC<=(REG[2] == REG[0])?PC+4+8*4:PC+4;
      10'h03e: data = 32'h00000000; // 004000f8: SLL, REG[0]<=REG[0]<<0;
      10'h03f: data = 32'h8fc40010; // 004000fc: LW, REG[4]<=RAM[REG[30]+16];
      10'h040: data = 32'h0c100174; // 00400100: JAL, PC<=0x00100174*4(=0x004005d0); REG[31]<=PC+4
      10'h041: data = 32'h00000000; // 00400104: SLL, REG[0]<=REG[0]<<0;
      10'h042: data = 32'h0c100066; // 00400108: JAL, PC<=0x00100066*4(=0x00400198); REG[31]<=PC+4
      10'h043: data = 32'h00000000; // 0040010c: SLL, REG[0]<=REG[0]<<0;
      10'h044: data = 32'h08100048; // 00400110: J, PC<=0x00100048*4(=0x00400120);
      10'h045: data = 32'h00000000; // 00400114: SLL, REG[0]<=REG[0]<<0;
      10'h046: data = 32'h0c10007c; // 00400118: JAL, PC<=0x0010007c*4(=0x004001f0); REG[31]<=PC+4
      10'h047: data = 32'h00000000; // 0040011c: SLL, REG[0]<=REG[0]<<0;
      10'h048: data = 32'h8fc20010; // 00400120: LW, REG[2]<=RAM[REG[30]+16];
      10'h049: data = 32'h00000000; // 00400124: SLL, REG[0]<=REG[0]<<0;
      10'h04a: data = 32'h24420001; // 00400128: ADDIU, REG[2]<=REG[2]+1(=0x00000001);
      10'h04b: data = 32'hafc20010; // 0040012c: SW, RAM[REG[30]+16]<=REG[2];
      10'h04c: data = 32'h8fc20010; // 00400130: LW, REG[2]<=RAM[REG[30]+16];
      10'h04d: data = 32'h00000000; // 00400134: SLL, REG[0]<=REG[0]<<0;
      10'h04e: data = 32'h2c420201; // 00400138: SLTIU, REG[2]<=(REG[2]<513(=0x00000201))?1:0;
      10'h04f: data = 32'h1440ffe9; // 0040013c: BNE, PC<=(REG[2] != REG[0])?PC+4+65513*4:PC+4;
      10'h050: data = 32'h00000000; // 00400140: SLL, REG[0]<=REG[0]<<0;
      10'h051: data = 32'h03c0e821; // 00400144: ADDU, REG[29]<=REG[30]+REG[0];
      10'h052: data = 32'h8fbf005c; // 00400148: LW, REG[31]<=RAM[REG[29]+92];
      10'h053: data = 32'h8fbe0058; // 0040014c: LW, REG[30]<=RAM[REG[29]+88];
      10'h054: data = 32'h27bd0060; // 00400150: ADDIU, REG[29]<=REG[29]+96(=0x00000060);
      10'h055: data = 32'h03e00008; // 00400154: JR, PC<=REG[31];
      10'h056: data = 32'h00000000; // 00400158: SLL, REG[0]<=REG[0]<<0;
      10'h057: data = 32'h27bdfff8; // 0040015c: ADDIU, REG[29]<=REG[29]+65528(=0x0000fff8);
      10'h058: data = 32'hafbe0000; // 00400160: SW, RAM[REG[29]+0]<=REG[30];
      10'h059: data = 32'h03a0f021; // 00400164: ADDU, REG[30]<=REG[29]+REG[0];
      10'h05a: data = 32'hafc40008; // 00400168: SW, RAM[REG[30]+8]<=REG[4];
      10'h05b: data = 32'h8fc20008; // 0040016c: LW, REG[2]<=RAM[REG[30]+8];
      10'h05c: data = 32'h00000000; // 00400170: SLL, REG[0]<=REG[0]<<0;
      10'h05d: data = 32'h8c420000; // 00400174: LW, REG[2]<=RAM[REG[2]+0];
      10'h05e: data = 32'h00000000; // 00400178: SLL, REG[0]<=REG[0]<<0;
      10'h05f: data = 32'h3842004e; // 0040017c: XORI
      10'h060: data = 32'h2c420001; // 00400180: SLTIU, REG[2]<=(REG[2]<1(=0x00000001))?1:0;
      10'h061: data = 32'h03c0e821; // 00400184: ADDU, REG[29]<=REG[30]+REG[0];
      10'h062: data = 32'h8fbe0000; // 00400188: LW, REG[30]<=RAM[REG[29]+0];
      10'h063: data = 32'h27bd0008; // 0040018c: ADDIU, REG[29]<=REG[29]+8(=0x00000008);
      10'h064: data = 32'h03e00008; // 00400190: JR, PC<=REG[31];
      10'h065: data = 32'h00000000; // 00400194: SLL, REG[0]<=REG[0]<<0;
      10'h066: data = 32'h27bdffe8; // 00400198: ADDIU, REG[29]<=REG[29]+65512(=0x0000ffe8);
      10'h067: data = 32'hafbf0014; // 0040019c: SW, RAM[REG[29]+20]<=REG[31];
      10'h068: data = 32'hafbe0010; // 004001a0: SW, RAM[REG[29]+16]<=REG[30];
      10'h069: data = 32'h03a0f021; // 004001a4: ADDU, REG[30]<=REG[29]+REG[0];
      10'h06a: data = 32'h24040008; // 004001a8: ADDIU, REG[4]<=REG[0]+8(=0x00000008);
      10'h06b: data = 32'h0c100241; // 004001ac: JAL, PC<=0x00100241*4(=0x00400904); REG[31]<=PC+4
      10'h06c: data = 32'h00000000; // 004001b0: SLL, REG[0]<=REG[0]<<0;
      10'h06d: data = 32'h24040004; // 004001b4: ADDIU, REG[4]<=REG[0]+4(=0x00000004);
      10'h06e: data = 32'h0c100241; // 004001b8: JAL, PC<=0x00100241*4(=0x00400904); REG[31]<=PC+4
      10'h06f: data = 32'h00000000; // 004001bc: SLL, REG[0]<=REG[0]<<0;
      10'h070: data = 32'h24040002; // 004001c0: ADDIU, REG[4]<=REG[0]+2(=0x00000002);
      10'h071: data = 32'h0c100241; // 004001c4: JAL, PC<=0x00100241*4(=0x00400904); REG[31]<=PC+4
      10'h072: data = 32'h00000000; // 004001c8: SLL, REG[0]<=REG[0]<<0;
      10'h073: data = 32'h24040001; // 004001cc: ADDIU, REG[4]<=REG[0]+1(=0x00000001);
      10'h074: data = 32'h0c100241; // 004001d0: JAL, PC<=0x00100241*4(=0x00400904); REG[31]<=PC+4
      10'h075: data = 32'h00000000; // 004001d4: SLL, REG[0]<=REG[0]<<0;
      10'h076: data = 32'h03c0e821; // 004001d8: ADDU, REG[29]<=REG[30]+REG[0];
      10'h077: data = 32'h8fbf0014; // 004001dc: LW, REG[31]<=RAM[REG[29]+20];
      10'h078: data = 32'h8fbe0010; // 004001e0: LW, REG[30]<=RAM[REG[29]+16];
      10'h079: data = 32'h27bd0018; // 004001e4: ADDIU, REG[29]<=REG[29]+24(=0x00000018);
      10'h07a: data = 32'h03e00008; // 004001e8: JR, PC<=REG[31];
      10'h07b: data = 32'h00000000; // 004001ec: SLL, REG[0]<=REG[0]<<0;
      10'h07c: data = 32'h27bdffe8; // 004001f0: ADDIU, REG[29]<=REG[29]+65512(=0x0000ffe8);
      10'h07d: data = 32'hafbf0014; // 004001f4: SW, RAM[REG[29]+20]<=REG[31];
      10'h07e: data = 32'hafbe0010; // 004001f8: SW, RAM[REG[29]+16]<=REG[30];
      10'h07f: data = 32'h03a0f021; // 004001fc: ADDU, REG[30]<=REG[29]+REG[0];
      10'h080: data = 32'h24040001; // 00400200: ADDIU, REG[4]<=REG[0]+1(=0x00000001);
      10'h081: data = 32'h0c100241; // 00400204: JAL, PC<=0x00100241*4(=0x00400904); REG[31]<=PC+4
      10'h082: data = 32'h00000000; // 00400208: SLL, REG[0]<=REG[0]<<0;
      10'h083: data = 32'h24040002; // 0040020c: ADDIU, REG[4]<=REG[0]+2(=0x00000002);
      10'h084: data = 32'h0c100241; // 00400210: JAL, PC<=0x00100241*4(=0x00400904); REG[31]<=PC+4
      10'h085: data = 32'h00000000; // 00400214: SLL, REG[0]<=REG[0]<<0;
      10'h086: data = 32'h24040004; // 00400218: ADDIU, REG[4]<=REG[0]+4(=0x00000004);
      10'h087: data = 32'h0c100241; // 0040021c: JAL, PC<=0x00100241*4(=0x00400904); REG[31]<=PC+4
      10'h088: data = 32'h00000000; // 00400220: SLL, REG[0]<=REG[0]<<0;
      10'h089: data = 32'h24040008; // 00400224: ADDIU, REG[4]<=REG[0]+8(=0x00000008);
      10'h08a: data = 32'h0c100241; // 00400228: JAL, PC<=0x00100241*4(=0x00400904); REG[31]<=PC+4
      10'h08b: data = 32'h00000000; // 0040022c: SLL, REG[0]<=REG[0]<<0;
      10'h08c: data = 32'h03c0e821; // 00400230: ADDU, REG[29]<=REG[30]+REG[0];
      10'h08d: data = 32'h8fbf0014; // 00400234: LW, REG[31]<=RAM[REG[29]+20];
      10'h08e: data = 32'h8fbe0010; // 00400238: LW, REG[30]<=RAM[REG[29]+16];
      10'h08f: data = 32'h27bd0018; // 0040023c: ADDIU, REG[29]<=REG[29]+24(=0x00000018);
      10'h090: data = 32'h03e00008; // 00400240: JR, PC<=REG[31];
      10'h091: data = 32'h00000000; // 00400244: SLL, REG[0]<=REG[0]<<0;
      10'h092: data = 32'h27bdfff8; // 00400248: ADDIU, REG[29]<=REG[29]+65528(=0x0000fff8);
      10'h093: data = 32'hafbe0000; // 0040024c: SW, RAM[REG[29]+0]<=REG[30];
      10'h094: data = 32'h03a0f021; // 00400250: ADDU, REG[30]<=REG[29]+REG[0];
      10'h095: data = 32'hafc40008; // 00400254: SW, RAM[REG[30]+8]<=REG[4];
      10'h096: data = 32'h24020308; // 00400258: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h097: data = 32'hac400000; // 0040025c: SW, RAM[REG[2]+0]<=REG[0];
      10'h098: data = 32'h2403030c; // 00400260: ADDIU, REG[3]<=REG[0]+780(=0x0000030c);
      10'h099: data = 32'h24020001; // 00400264: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h09a: data = 32'hac620000; // 00400268: SW, RAM[REG[3]+0]<=REG[2];
      10'h09b: data = 32'h24030308; // 0040026c: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h09c: data = 32'h24020001; // 00400270: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h09d: data = 32'hac620000; // 00400274: SW, RAM[REG[3]+0]<=REG[2];
      10'h09e: data = 32'h24020308; // 00400278: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h09f: data = 32'hac400000; // 0040027c: SW, RAM[REG[2]+0]<=REG[0];
      10'h0a0: data = 32'h24030308; // 00400280: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h0a1: data = 32'h24020001; // 00400284: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h0a2: data = 32'hac620000; // 00400288: SW, RAM[REG[3]+0]<=REG[2];
      10'h0a3: data = 32'h081000aa; // 0040028c: J, PC<=0x001000aa*4(=0x004002a8);
      10'h0a4: data = 32'h00000000; // 00400290: SLL, REG[0]<=REG[0]<<0;
      10'h0a5: data = 32'h24020308; // 00400294: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h0a6: data = 32'hac400000; // 00400298: SW, RAM[REG[2]+0]<=REG[0];
      10'h0a7: data = 32'h24030308; // 0040029c: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h0a8: data = 32'h24020001; // 004002a0: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h0a9: data = 32'hac620000; // 004002a4: SW, RAM[REG[3]+0]<=REG[2];
      10'h0aa: data = 32'h24020310; // 004002a8: ADDIU, REG[2]<=REG[0]+784(=0x00000310);
      10'h0ab: data = 32'h8c430000; // 004002ac: LW, REG[3]<=RAM[REG[2]+0];
      10'h0ac: data = 32'h2402ffff; // 004002b0: ADDIU, REG[2]<=REG[0]+65535(=0x0000ffff);
      10'h0ad: data = 32'h1062fff7; // 004002b4: BEQ, PC<=(REG[3] == REG[2])?PC+4+65527*4:PC+4;
      10'h0ae: data = 32'h00000000; // 004002b8: SLL, REG[0]<=REG[0]<<0;
      10'h0af: data = 32'h08100158; // 004002bc: J, PC<=0x00100158*4(=0x00400560);
      10'h0b0: data = 32'h00000000; // 004002c0: SLL, REG[0]<=REG[0]<<0;
      10'h0b1: data = 32'h8fc20008; // 004002c4: LW, REG[2]<=RAM[REG[30]+8];
      10'h0b2: data = 32'h00000000; // 004002c8: SLL, REG[0]<=REG[0]<<0;
      10'h0b3: data = 32'h8c420000; // 004002cc: LW, REG[2]<=RAM[REG[2]+0];
      10'h0b4: data = 32'h00000000; // 004002d0: SLL, REG[0]<=REG[0]<<0;
      10'h0b5: data = 32'h10400012; // 004002d4: BEQ, PC<=(REG[2] == REG[0])?PC+4+18*4:PC+4;
      10'h0b6: data = 32'h00000000; // 004002d8: SLL, REG[0]<=REG[0]<<0;
      10'h0b7: data = 32'h8fc20008; // 004002dc: LW, REG[2]<=RAM[REG[30]+8];
      10'h0b8: data = 32'h00000000; // 004002e0: SLL, REG[0]<=REG[0]<<0;
      10'h0b9: data = 32'h8c420000; // 004002e4: LW, REG[2]<=RAM[REG[2]+0];
      10'h0ba: data = 32'h00000000; // 004002e8: SLL, REG[0]<=REG[0]<<0;
      10'h0bb: data = 32'h2c42001b; // 004002ec: SLTIU, REG[2]<=(REG[2]<27(=0x0000001b))?1:0;
      10'h0bc: data = 32'h1040000b; // 004002f0: BEQ, PC<=(REG[2] == REG[0])?PC+4+11*4:PC+4;
      10'h0bd: data = 32'h00000000; // 004002f4: SLL, REG[0]<=REG[0]<<0;
      10'h0be: data = 32'h8fc20008; // 004002f8: LW, REG[2]<=RAM[REG[30]+8];
      10'h0bf: data = 32'h00000000; // 004002fc: SLL, REG[0]<=REG[0]<<0;
      10'h0c0: data = 32'h8c420000; // 00400300: LW, REG[2]<=RAM[REG[2]+0];
      10'h0c1: data = 32'h00000000; // 00400304: SLL, REG[0]<=REG[0]<<0;
      10'h0c2: data = 32'h24430040; // 00400308: ADDIU, REG[3]<=REG[2]+64(=0x00000040);
      10'h0c3: data = 32'h8fc20008; // 0040030c: LW, REG[2]<=RAM[REG[30]+8];
      10'h0c4: data = 32'h00000000; // 00400310: SLL, REG[0]<=REG[0]<<0;
      10'h0c5: data = 32'hac430000; // 00400314: SW, RAM[REG[2]+0]<=REG[3];
      10'h0c6: data = 32'h0810014f; // 00400318: J, PC<=0x0010014f*4(=0x0040053c);
      10'h0c7: data = 32'h00000000; // 0040031c: SLL, REG[0]<=REG[0]<<0;
      10'h0c8: data = 32'h8fc20008; // 00400320: LW, REG[2]<=RAM[REG[30]+8];
      10'h0c9: data = 32'h00000000; // 00400324: SLL, REG[0]<=REG[0]<<0;
      10'h0ca: data = 32'h8c420000; // 00400328: LW, REG[2]<=RAM[REG[2]+0];
      10'h0cb: data = 32'h00000000; // 0040032c: SLL, REG[0]<=REG[0]<<0;
      10'h0cc: data = 32'h2c420030; // 00400330: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h0cd: data = 32'h14400010; // 00400334: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h0ce: data = 32'h00000000; // 00400338: SLL, REG[0]<=REG[0]<<0;
      10'h0cf: data = 32'h8fc20008; // 0040033c: LW, REG[2]<=RAM[REG[30]+8];
      10'h0d0: data = 32'h00000000; // 00400340: SLL, REG[0]<=REG[0]<<0;
      10'h0d1: data = 32'h8c420000; // 00400344: LW, REG[2]<=RAM[REG[2]+0];
      10'h0d2: data = 32'h00000000; // 00400348: SLL, REG[0]<=REG[0]<<0;
      10'h0d3: data = 32'h2c42003a; // 0040034c: SLTIU, REG[2]<=(REG[2]<58(=0x0000003a))?1:0;
      10'h0d4: data = 32'h10400009; // 00400350: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h0d5: data = 32'h00000000; // 00400354: SLL, REG[0]<=REG[0]<<0;
      10'h0d6: data = 32'h8fc20008; // 00400358: LW, REG[2]<=RAM[REG[30]+8];
      10'h0d7: data = 32'h00000000; // 0040035c: SLL, REG[0]<=REG[0]<<0;
      10'h0d8: data = 32'h8c430000; // 00400360: LW, REG[3]<=RAM[REG[2]+0];
      10'h0d9: data = 32'h8fc20008; // 00400364: LW, REG[2]<=RAM[REG[30]+8];
      10'h0da: data = 32'h00000000; // 00400368: SLL, REG[0]<=REG[0]<<0;
      10'h0db: data = 32'hac430000; // 0040036c: SW, RAM[REG[2]+0]<=REG[3];
      10'h0dc: data = 32'h0810014f; // 00400370: J, PC<=0x0010014f*4(=0x0040053c);
      10'h0dd: data = 32'h00000000; // 00400374: SLL, REG[0]<=REG[0]<<0;
      10'h0de: data = 32'h8fc20008; // 00400378: LW, REG[2]<=RAM[REG[30]+8];
      10'h0df: data = 32'h00000000; // 0040037c: SLL, REG[0]<=REG[0]<<0;
      10'h0e0: data = 32'h8c420000; // 00400380: LW, REG[2]<=RAM[REG[2]+0];
      10'h0e1: data = 32'h00000000; // 00400384: SLL, REG[0]<=REG[0]<<0;
      10'h0e2: data = 32'h14400006; // 00400388: BNE, PC<=(REG[2] != REG[0])?PC+4+6*4:PC+4;
      10'h0e3: data = 32'h00000000; // 0040038c: SLL, REG[0]<=REG[0]<<0;
      10'h0e4: data = 32'h8fc30008; // 00400390: LW, REG[3]<=RAM[REG[30]+8];
      10'h0e5: data = 32'h24020040; // 00400394: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h0e6: data = 32'hac620000; // 00400398: SW, RAM[REG[3]+0]<=REG[2];
      10'h0e7: data = 32'h0810014f; // 0040039c: J, PC<=0x0010014f*4(=0x0040053c);
      10'h0e8: data = 32'h00000000; // 004003a0: SLL, REG[0]<=REG[0]<<0;
      10'h0e9: data = 32'h8fc20008; // 004003a4: LW, REG[2]<=RAM[REG[30]+8];
      10'h0ea: data = 32'h00000000; // 004003a8: SLL, REG[0]<=REG[0]<<0;
      10'h0eb: data = 32'h8c430000; // 004003ac: LW, REG[3]<=RAM[REG[2]+0];
      10'h0ec: data = 32'h2402001b; // 004003b0: ADDIU, REG[2]<=REG[0]+27(=0x0000001b);
      10'h0ed: data = 32'h14620006; // 004003b4: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0ee: data = 32'h00000000; // 004003b8: SLL, REG[0]<=REG[0]<<0;
      10'h0ef: data = 32'h8fc30008; // 004003bc: LW, REG[3]<=RAM[REG[30]+8];
      10'h0f0: data = 32'h2402005b; // 004003c0: ADDIU, REG[2]<=REG[0]+91(=0x0000005b);
      10'h0f1: data = 32'hac620000; // 004003c4: SW, RAM[REG[3]+0]<=REG[2];
      10'h0f2: data = 32'h0810014f; // 004003c8: J, PC<=0x0010014f*4(=0x0040053c);
      10'h0f3: data = 32'h00000000; // 004003cc: SLL, REG[0]<=REG[0]<<0;
      10'h0f4: data = 32'h8fc20008; // 004003d0: LW, REG[2]<=RAM[REG[30]+8];
      10'h0f5: data = 32'h00000000; // 004003d4: SLL, REG[0]<=REG[0]<<0;
      10'h0f6: data = 32'h8c430000; // 004003d8: LW, REG[3]<=RAM[REG[2]+0];
      10'h0f7: data = 32'h2402001d; // 004003dc: ADDIU, REG[2]<=REG[0]+29(=0x0000001d);
      10'h0f8: data = 32'h14620006; // 004003e0: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h0f9: data = 32'h00000000; // 004003e4: SLL, REG[0]<=REG[0]<<0;
      10'h0fa: data = 32'h8fc30008; // 004003e8: LW, REG[3]<=RAM[REG[30]+8];
      10'h0fb: data = 32'h2402005d; // 004003ec: ADDIU, REG[2]<=REG[0]+93(=0x0000005d);
      10'h0fc: data = 32'hac620000; // 004003f0: SW, RAM[REG[3]+0]<=REG[2];
      10'h0fd: data = 32'h0810014f; // 004003f4: J, PC<=0x0010014f*4(=0x0040053c);
      10'h0fe: data = 32'h00000000; // 004003f8: SLL, REG[0]<=REG[0]<<0;
      10'h0ff: data = 32'h8fc20008; // 004003fc: LW, REG[2]<=RAM[REG[30]+8];
      10'h100: data = 32'h00000000; // 00400400: SLL, REG[0]<=REG[0]<<0;
      10'h101: data = 32'h8c420000; // 00400404: LW, REG[2]<=RAM[REG[2]+0];
      10'h102: data = 32'h00000000; // 00400408: SLL, REG[0]<=REG[0]<<0;
      10'h103: data = 32'h2c420020; // 0040040c: SLTIU, REG[2]<=(REG[2]<32(=0x00000020))?1:0;
      10'h104: data = 32'h14400010; // 00400410: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h105: data = 32'h00000000; // 00400414: SLL, REG[0]<=REG[0]<<0;
      10'h106: data = 32'h8fc20008; // 00400418: LW, REG[2]<=RAM[REG[30]+8];
      10'h107: data = 32'h00000000; // 0040041c: SLL, REG[0]<=REG[0]<<0;
      10'h108: data = 32'h8c420000; // 00400420: LW, REG[2]<=RAM[REG[2]+0];
      10'h109: data = 32'h00000000; // 00400424: SLL, REG[0]<=REG[0]<<0;
      10'h10a: data = 32'h2c420030; // 00400428: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h10b: data = 32'h10400009; // 0040042c: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h10c: data = 32'h00000000; // 00400430: SLL, REG[0]<=REG[0]<<0;
      10'h10d: data = 32'h8fc20008; // 00400434: LW, REG[2]<=RAM[REG[30]+8];
      10'h10e: data = 32'h00000000; // 00400438: SLL, REG[0]<=REG[0]<<0;
      10'h10f: data = 32'h8c430000; // 0040043c: LW, REG[3]<=RAM[REG[2]+0];
      10'h110: data = 32'h8fc20008; // 00400440: LW, REG[2]<=RAM[REG[30]+8];
      10'h111: data = 32'h00000000; // 00400444: SLL, REG[0]<=REG[0]<<0;
      10'h112: data = 32'hac430000; // 00400448: SW, RAM[REG[2]+0]<=REG[3];
      10'h113: data = 32'h0810014f; // 0040044c: J, PC<=0x0010014f*4(=0x0040053c);
      10'h114: data = 32'h00000000; // 00400450: SLL, REG[0]<=REG[0]<<0;
      10'h115: data = 32'h8fc20008; // 00400454: LW, REG[2]<=RAM[REG[30]+8];
      10'h116: data = 32'h00000000; // 00400458: SLL, REG[0]<=REG[0]<<0;
      10'h117: data = 32'h8c430000; // 0040045c: LW, REG[3]<=RAM[REG[2]+0];
      10'h118: data = 32'h2402003a; // 00400460: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h119: data = 32'h14620006; // 00400464: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h11a: data = 32'h00000000; // 00400468: SLL, REG[0]<=REG[0]<<0;
      10'h11b: data = 32'h8fc30008; // 0040046c: LW, REG[3]<=RAM[REG[30]+8];
      10'h11c: data = 32'h2402003f; // 00400470: ADDIU, REG[2]<=REG[0]+63(=0x0000003f);
      10'h11d: data = 32'hac620000; // 00400474: SW, RAM[REG[3]+0]<=REG[2];
      10'h11e: data = 32'h0810014f; // 00400478: J, PC<=0x0010014f*4(=0x0040053c);
      10'h11f: data = 32'h00000000; // 0040047c: SLL, REG[0]<=REG[0]<<0;
      10'h120: data = 32'h8fc20008; // 00400480: LW, REG[2]<=RAM[REG[30]+8];
      10'h121: data = 32'h00000000; // 00400484: SLL, REG[0]<=REG[0]<<0;
      10'h122: data = 32'h8c430000; // 00400488: LW, REG[3]<=RAM[REG[2]+0];
      10'h123: data = 32'h2402003b; // 0040048c: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h124: data = 32'h14620006; // 00400490: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h125: data = 32'h00000000; // 00400494: SLL, REG[0]<=REG[0]<<0;
      10'h126: data = 32'h8fc30008; // 00400498: LW, REG[3]<=RAM[REG[30]+8];
      10'h127: data = 32'h2402003d; // 0040049c: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h128: data = 32'hac620000; // 004004a0: SW, RAM[REG[3]+0]<=REG[2];
      10'h129: data = 32'h0810014f; // 004004a4: J, PC<=0x0010014f*4(=0x0040053c);
      10'h12a: data = 32'h00000000; // 004004a8: SLL, REG[0]<=REG[0]<<0;
      10'h12b: data = 32'h8fc20008; // 004004ac: LW, REG[2]<=RAM[REG[30]+8];
      10'h12c: data = 32'h00000000; // 004004b0: SLL, REG[0]<=REG[0]<<0;
      10'h12d: data = 32'h8c430000; // 004004b4: LW, REG[3]<=RAM[REG[2]+0];
      10'h12e: data = 32'h2402003c; // 004004b8: ADDIU, REG[2]<=REG[0]+60(=0x0000003c);
      10'h12f: data = 32'h14620006; // 004004bc: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h130: data = 32'h00000000; // 004004c0: SLL, REG[0]<=REG[0]<<0;
      10'h131: data = 32'h8fc30008; // 004004c4: LW, REG[3]<=RAM[REG[30]+8];
      10'h132: data = 32'h2402003b; // 004004c8: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h133: data = 32'hac620000; // 004004cc: SW, RAM[REG[3]+0]<=REG[2];
      10'h134: data = 32'h0810014f; // 004004d0: J, PC<=0x0010014f*4(=0x0040053c);
      10'h135: data = 32'h00000000; // 004004d4: SLL, REG[0]<=REG[0]<<0;
      10'h136: data = 32'h8fc20008; // 004004d8: LW, REG[2]<=RAM[REG[30]+8];
      10'h137: data = 32'h00000000; // 004004dc: SLL, REG[0]<=REG[0]<<0;
      10'h138: data = 32'h8c430000; // 004004e0: LW, REG[3]<=RAM[REG[2]+0];
      10'h139: data = 32'h2402003d; // 004004e4: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h13a: data = 32'h14620006; // 004004e8: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h13b: data = 32'h00000000; // 004004ec: SLL, REG[0]<=REG[0]<<0;
      10'h13c: data = 32'h8fc30008; // 004004f0: LW, REG[3]<=RAM[REG[30]+8];
      10'h13d: data = 32'h2402003a; // 004004f4: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h13e: data = 32'hac620000; // 004004f8: SW, RAM[REG[3]+0]<=REG[2];
      10'h13f: data = 32'h0810014f; // 004004fc: J, PC<=0x0010014f*4(=0x0040053c);
      10'h140: data = 32'h00000000; // 00400500: SLL, REG[0]<=REG[0]<<0;
      10'h141: data = 32'h8fc20008; // 00400504: LW, REG[2]<=RAM[REG[30]+8];
      10'h142: data = 32'h00000000; // 00400508: SLL, REG[0]<=REG[0]<<0;
      10'h143: data = 32'h8c430000; // 0040050c: LW, REG[3]<=RAM[REG[2]+0];
      10'h144: data = 32'h2402003e; // 00400510: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h145: data = 32'h14620006; // 00400514: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h146: data = 32'h00000000; // 00400518: SLL, REG[0]<=REG[0]<<0;
      10'h147: data = 32'h8fc30008; // 0040051c: LW, REG[3]<=RAM[REG[30]+8];
      10'h148: data = 32'h2402000a; // 00400520: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h149: data = 32'hac620000; // 00400524: SW, RAM[REG[3]+0]<=REG[2];
      10'h14a: data = 32'h0810014f; // 00400528: J, PC<=0x0010014f*4(=0x0040053c);
      10'h14b: data = 32'h00000000; // 0040052c: SLL, REG[0]<=REG[0]<<0;
      10'h14c: data = 32'h8fc30008; // 00400530: LW, REG[3]<=RAM[REG[30]+8];
      10'h14d: data = 32'h24020040; // 00400534: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h14e: data = 32'hac620000; // 00400538: SW, RAM[REG[3]+0]<=REG[2];
      10'h14f: data = 32'h24020308; // 0040053c: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h150: data = 32'hac400000; // 00400540: SW, RAM[REG[2]+0]<=REG[0];
      10'h151: data = 32'h24030308; // 00400544: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h152: data = 32'h24020001; // 00400548: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h153: data = 32'hac620000; // 0040054c: SW, RAM[REG[3]+0]<=REG[2];
      10'h154: data = 32'h8fc20008; // 00400550: LW, REG[2]<=RAM[REG[30]+8];
      10'h155: data = 32'h00000000; // 00400554: SLL, REG[0]<=REG[0]<<0;
      10'h156: data = 32'h24420004; // 00400558: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h157: data = 32'hafc20008; // 0040055c: SW, RAM[REG[30]+8]<=REG[2];
      10'h158: data = 32'h24020310; // 00400560: ADDIU, REG[2]<=REG[0]+784(=0x00000310);
      10'h159: data = 32'h8c430000; // 00400564: LW, REG[3]<=RAM[REG[2]+0];
      10'h15a: data = 32'h8fc20008; // 00400568: LW, REG[2]<=RAM[REG[30]+8];
      10'h15b: data = 32'h00000000; // 0040056c: SLL, REG[0]<=REG[0]<<0;
      10'h15c: data = 32'hac430000; // 00400570: SW, RAM[REG[2]+0]<=REG[3];
      10'h15d: data = 32'h8fc20008; // 00400574: LW, REG[2]<=RAM[REG[30]+8];
      10'h15e: data = 32'h00000000; // 00400578: SLL, REG[0]<=REG[0]<<0;
      10'h15f: data = 32'h8c430000; // 0040057c: LW, REG[3]<=RAM[REG[2]+0];
      10'h160: data = 32'h2402003e; // 00400580: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h161: data = 32'h1462ff4f; // 00400584: BNE, PC<=(REG[3] != REG[2])?PC+4+65359*4:PC+4;
      10'h162: data = 32'h00000000; // 00400588: SLL, REG[0]<=REG[0]<<0;
      10'h163: data = 32'h8fc20008; // 0040058c: LW, REG[2]<=RAM[REG[30]+8];
      10'h164: data = 32'h00000000; // 00400590: SLL, REG[0]<=REG[0]<<0;
      10'h165: data = 32'hac400000; // 00400594: SW, RAM[REG[2]+0]<=REG[0];
      10'h166: data = 32'h24020308; // 00400598: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h167: data = 32'hac400000; // 0040059c: SW, RAM[REG[2]+0]<=REG[0];
      10'h168: data = 32'h2402030c; // 004005a0: ADDIU, REG[2]<=REG[0]+780(=0x0000030c);
      10'h169: data = 32'hac400000; // 004005a4: SW, RAM[REG[2]+0]<=REG[0];
      10'h16a: data = 32'h24030308; // 004005a8: ADDIU, REG[3]<=REG[0]+776(=0x00000308);
      10'h16b: data = 32'h24020001; // 004005ac: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h16c: data = 32'hac620000; // 004005b0: SW, RAM[REG[3]+0]<=REG[2];
      10'h16d: data = 32'h24020308; // 004005b4: ADDIU, REG[2]<=REG[0]+776(=0x00000308);
      10'h16e: data = 32'hac400000; // 004005b8: SW, RAM[REG[2]+0]<=REG[0];
      10'h16f: data = 32'h03c0e821; // 004005bc: ADDU, REG[29]<=REG[30]+REG[0];
      10'h170: data = 32'h8fbe0000; // 004005c0: LW, REG[30]<=RAM[REG[29]+0];
      10'h171: data = 32'h27bd0008; // 004005c4: ADDIU, REG[29]<=REG[29]+8(=0x00000008);
      10'h172: data = 32'h03e00008; // 004005c8: JR, PC<=REG[31];
      10'h173: data = 32'h00000000; // 004005cc: SLL, REG[0]<=REG[0]<<0;
      10'h174: data = 32'h27bdfff8; // 004005d0: ADDIU, REG[29]<=REG[29]+65528(=0x0000fff8);
      10'h175: data = 32'hafbe0000; // 004005d4: SW, RAM[REG[29]+0]<=REG[30];
      10'h176: data = 32'h03a0f021; // 004005d8: ADDU, REG[30]<=REG[29]+REG[0];
      10'h177: data = 32'hafc40008; // 004005dc: SW, RAM[REG[30]+8]<=REG[4];
      10'h178: data = 32'h08100236; // 004005e0: J, PC<=0x00100236*4(=0x004008d8);
      10'h179: data = 32'h00000000; // 004005e4: SLL, REG[0]<=REG[0]<<0;
      10'h17a: data = 32'h24020300; // 004005e8: ADDIU, REG[2]<=REG[0]+768(=0x00000300);
      10'h17b: data = 32'hac400000; // 004005ec: SW, RAM[REG[2]+0]<=REG[0];
      10'h17c: data = 32'h8fc20008; // 004005f0: LW, REG[2]<=RAM[REG[30]+8];
      10'h17d: data = 32'h00000000; // 004005f4: SLL, REG[0]<=REG[0]<<0;
      10'h17e: data = 32'h8c420000; // 004005f8: LW, REG[2]<=RAM[REG[2]+0];
      10'h17f: data = 32'h00000000; // 004005fc: SLL, REG[0]<=REG[0]<<0;
      10'h180: data = 32'h2c420041; // 00400600: SLTIU, REG[2]<=(REG[2]<65(=0x00000041))?1:0;
      10'h181: data = 32'h14400011; // 00400604: BNE, PC<=(REG[2] != REG[0])?PC+4+17*4:PC+4;
      10'h182: data = 32'h00000000; // 00400608: SLL, REG[0]<=REG[0]<<0;
      10'h183: data = 32'h8fc20008; // 0040060c: LW, REG[2]<=RAM[REG[30]+8];
      10'h184: data = 32'h00000000; // 00400610: SLL, REG[0]<=REG[0]<<0;
      10'h185: data = 32'h8c420000; // 00400614: LW, REG[2]<=RAM[REG[2]+0];
      10'h186: data = 32'h00000000; // 00400618: SLL, REG[0]<=REG[0]<<0;
      10'h187: data = 32'h2c42005b; // 0040061c: SLTIU, REG[2]<=(REG[2]<91(=0x0000005b))?1:0;
      10'h188: data = 32'h1040000a; // 00400620: BEQ, PC<=(REG[2] == REG[0])?PC+4+10*4:PC+4;
      10'h189: data = 32'h00000000; // 00400624: SLL, REG[0]<=REG[0]<<0;
      10'h18a: data = 32'h24030304; // 00400628: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h18b: data = 32'h8fc20008; // 0040062c: LW, REG[2]<=RAM[REG[30]+8];
      10'h18c: data = 32'h00000000; // 00400630: SLL, REG[0]<=REG[0]<<0;
      10'h18d: data = 32'h8c420000; // 00400634: LW, REG[2]<=RAM[REG[2]+0];
      10'h18e: data = 32'h00000000; // 00400638: SLL, REG[0]<=REG[0]<<0;
      10'h18f: data = 32'h2442ffc0; // 0040063c: ADDIU, REG[2]<=REG[2]+65472(=0x0000ffc0);
      10'h190: data = 32'hac620000; // 00400640: SW, RAM[REG[3]+0]<=REG[2];
      10'h191: data = 32'h0810022f; // 00400644: J, PC<=0x0010022f*4(=0x004008bc);
      10'h192: data = 32'h00000000; // 00400648: SLL, REG[0]<=REG[0]<<0;
      10'h193: data = 32'h8fc20008; // 0040064c: LW, REG[2]<=RAM[REG[30]+8];
      10'h194: data = 32'h00000000; // 00400650: SLL, REG[0]<=REG[0]<<0;
      10'h195: data = 32'h8c420000; // 00400654: LW, REG[2]<=RAM[REG[2]+0];
      10'h196: data = 32'h00000000; // 00400658: SLL, REG[0]<=REG[0]<<0;
      10'h197: data = 32'h2c420061; // 0040065c: SLTIU, REG[2]<=(REG[2]<97(=0x00000061))?1:0;
      10'h198: data = 32'h14400011; // 00400660: BNE, PC<=(REG[2] != REG[0])?PC+4+17*4:PC+4;
      10'h199: data = 32'h00000000; // 00400664: SLL, REG[0]<=REG[0]<<0;
      10'h19a: data = 32'h8fc20008; // 00400668: LW, REG[2]<=RAM[REG[30]+8];
      10'h19b: data = 32'h00000000; // 0040066c: SLL, REG[0]<=REG[0]<<0;
      10'h19c: data = 32'h8c420000; // 00400670: LW, REG[2]<=RAM[REG[2]+0];
      10'h19d: data = 32'h00000000; // 00400674: SLL, REG[0]<=REG[0]<<0;
      10'h19e: data = 32'h2c42007b; // 00400678: SLTIU, REG[2]<=(REG[2]<123(=0x0000007b))?1:0;
      10'h19f: data = 32'h1040000a; // 0040067c: BEQ, PC<=(REG[2] == REG[0])?PC+4+10*4:PC+4;
      10'h1a0: data = 32'h00000000; // 00400680: SLL, REG[0]<=REG[0]<<0;
      10'h1a1: data = 32'h24030304; // 00400684: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h1a2: data = 32'h8fc20008; // 00400688: LW, REG[2]<=RAM[REG[30]+8];
      10'h1a3: data = 32'h00000000; // 0040068c: SLL, REG[0]<=REG[0]<<0;
      10'h1a4: data = 32'h8c420000; // 00400690: LW, REG[2]<=RAM[REG[2]+0];
      10'h1a5: data = 32'h00000000; // 00400694: SLL, REG[0]<=REG[0]<<0;
      10'h1a6: data = 32'h2442ffa0; // 00400698: ADDIU, REG[2]<=REG[2]+65440(=0x0000ffa0);
      10'h1a7: data = 32'hac620000; // 0040069c: SW, RAM[REG[3]+0]<=REG[2];
      10'h1a8: data = 32'h0810022f; // 004006a0: J, PC<=0x0010022f*4(=0x004008bc);
      10'h1a9: data = 32'h00000000; // 004006a4: SLL, REG[0]<=REG[0]<<0;
      10'h1aa: data = 32'h8fc20008; // 004006a8: LW, REG[2]<=RAM[REG[30]+8];
      10'h1ab: data = 32'h00000000; // 004006ac: SLL, REG[0]<=REG[0]<<0;
      10'h1ac: data = 32'h8c420000; // 004006b0: LW, REG[2]<=RAM[REG[2]+0];
      10'h1ad: data = 32'h00000000; // 004006b4: SLL, REG[0]<=REG[0]<<0;
      10'h1ae: data = 32'h2c420030; // 004006b8: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h1af: data = 32'h14400010; // 004006bc: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h1b0: data = 32'h00000000; // 004006c0: SLL, REG[0]<=REG[0]<<0;
      10'h1b1: data = 32'h8fc20008; // 004006c4: LW, REG[2]<=RAM[REG[30]+8];
      10'h1b2: data = 32'h00000000; // 004006c8: SLL, REG[0]<=REG[0]<<0;
      10'h1b3: data = 32'h8c420000; // 004006cc: LW, REG[2]<=RAM[REG[2]+0];
      10'h1b4: data = 32'h00000000; // 004006d0: SLL, REG[0]<=REG[0]<<0;
      10'h1b5: data = 32'h2c42003a; // 004006d4: SLTIU, REG[2]<=(REG[2]<58(=0x0000003a))?1:0;
      10'h1b6: data = 32'h10400009; // 004006d8: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h1b7: data = 32'h00000000; // 004006dc: SLL, REG[0]<=REG[0]<<0;
      10'h1b8: data = 32'h24020304; // 004006e0: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h1b9: data = 32'h8fc30008; // 004006e4: LW, REG[3]<=RAM[REG[30]+8];
      10'h1ba: data = 32'h00000000; // 004006e8: SLL, REG[0]<=REG[0]<<0;
      10'h1bb: data = 32'h8c630000; // 004006ec: LW, REG[3]<=RAM[REG[3]+0];
      10'h1bc: data = 32'h00000000; // 004006f0: SLL, REG[0]<=REG[0]<<0;
      10'h1bd: data = 32'hac430000; // 004006f4: SW, RAM[REG[2]+0]<=REG[3];
      10'h1be: data = 32'h0810022f; // 004006f8: J, PC<=0x0010022f*4(=0x004008bc);
      10'h1bf: data = 32'h00000000; // 004006fc: SLL, REG[0]<=REG[0]<<0;
      10'h1c0: data = 32'h8fc20008; // 00400700: LW, REG[2]<=RAM[REG[30]+8];
      10'h1c1: data = 32'h00000000; // 00400704: SLL, REG[0]<=REG[0]<<0;
      10'h1c2: data = 32'h8c430000; // 00400708: LW, REG[3]<=RAM[REG[2]+0];
      10'h1c3: data = 32'h24020040; // 0040070c: ADDIU, REG[2]<=REG[0]+64(=0x00000040);
      10'h1c4: data = 32'h14620005; // 00400710: BNE, PC<=(REG[3] != REG[2])?PC+4+5*4:PC+4;
      10'h1c5: data = 32'h00000000; // 00400714: SLL, REG[0]<=REG[0]<<0;
      10'h1c6: data = 32'h24020304; // 00400718: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h1c7: data = 32'hac400000; // 0040071c: SW, RAM[REG[2]+0]<=REG[0];
      10'h1c8: data = 32'h0810022f; // 00400720: J, PC<=0x0010022f*4(=0x004008bc);
      10'h1c9: data = 32'h00000000; // 00400724: SLL, REG[0]<=REG[0]<<0;
      10'h1ca: data = 32'h8fc20008; // 00400728: LW, REG[2]<=RAM[REG[30]+8];
      10'h1cb: data = 32'h00000000; // 0040072c: SLL, REG[0]<=REG[0]<<0;
      10'h1cc: data = 32'h8c430000; // 00400730: LW, REG[3]<=RAM[REG[2]+0];
      10'h1cd: data = 32'h2402005b; // 00400734: ADDIU, REG[2]<=REG[0]+91(=0x0000005b);
      10'h1ce: data = 32'h14620006; // 00400738: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h1cf: data = 32'h00000000; // 0040073c: SLL, REG[0]<=REG[0]<<0;
      10'h1d0: data = 32'h24030304; // 00400740: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h1d1: data = 32'h2402001b; // 00400744: ADDIU, REG[2]<=REG[0]+27(=0x0000001b);
      10'h1d2: data = 32'hac620000; // 00400748: SW, RAM[REG[3]+0]<=REG[2];
      10'h1d3: data = 32'h0810022f; // 0040074c: J, PC<=0x0010022f*4(=0x004008bc);
      10'h1d4: data = 32'h00000000; // 00400750: SLL, REG[0]<=REG[0]<<0;
      10'h1d5: data = 32'h8fc20008; // 00400754: LW, REG[2]<=RAM[REG[30]+8];
      10'h1d6: data = 32'h00000000; // 00400758: SLL, REG[0]<=REG[0]<<0;
      10'h1d7: data = 32'h8c430000; // 0040075c: LW, REG[3]<=RAM[REG[2]+0];
      10'h1d8: data = 32'h2402005d; // 00400760: ADDIU, REG[2]<=REG[0]+93(=0x0000005d);
      10'h1d9: data = 32'h14620006; // 00400764: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h1da: data = 32'h00000000; // 00400768: SLL, REG[0]<=REG[0]<<0;
      10'h1db: data = 32'h24030304; // 0040076c: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h1dc: data = 32'h2402001d; // 00400770: ADDIU, REG[2]<=REG[0]+29(=0x0000001d);
      10'h1dd: data = 32'hac620000; // 00400774: SW, RAM[REG[3]+0]<=REG[2];
      10'h1de: data = 32'h0810022f; // 00400778: J, PC<=0x0010022f*4(=0x004008bc);
      10'h1df: data = 32'h00000000; // 0040077c: SLL, REG[0]<=REG[0]<<0;
      10'h1e0: data = 32'h8fc20008; // 00400780: LW, REG[2]<=RAM[REG[30]+8];
      10'h1e1: data = 32'h00000000; // 00400784: SLL, REG[0]<=REG[0]<<0;
      10'h1e2: data = 32'h8c420000; // 00400788: LW, REG[2]<=RAM[REG[2]+0];
      10'h1e3: data = 32'h00000000; // 0040078c: SLL, REG[0]<=REG[0]<<0;
      10'h1e4: data = 32'h2c420020; // 00400790: SLTIU, REG[2]<=(REG[2]<32(=0x00000020))?1:0;
      10'h1e5: data = 32'h14400010; // 00400794: BNE, PC<=(REG[2] != REG[0])?PC+4+16*4:PC+4;
      10'h1e6: data = 32'h00000000; // 00400798: SLL, REG[0]<=REG[0]<<0;
      10'h1e7: data = 32'h8fc20008; // 0040079c: LW, REG[2]<=RAM[REG[30]+8];
      10'h1e8: data = 32'h00000000; // 004007a0: SLL, REG[0]<=REG[0]<<0;
      10'h1e9: data = 32'h8c420000; // 004007a4: LW, REG[2]<=RAM[REG[2]+0];
      10'h1ea: data = 32'h00000000; // 004007a8: SLL, REG[0]<=REG[0]<<0;
      10'h1eb: data = 32'h2c420030; // 004007ac: SLTIU, REG[2]<=(REG[2]<48(=0x00000030))?1:0;
      10'h1ec: data = 32'h10400009; // 004007b0: BEQ, PC<=(REG[2] == REG[0])?PC+4+9*4:PC+4;
      10'h1ed: data = 32'h00000000; // 004007b4: SLL, REG[0]<=REG[0]<<0;
      10'h1ee: data = 32'h24020304; // 004007b8: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h1ef: data = 32'h8fc30008; // 004007bc: LW, REG[3]<=RAM[REG[30]+8];
      10'h1f0: data = 32'h00000000; // 004007c0: SLL, REG[0]<=REG[0]<<0;
      10'h1f1: data = 32'h8c630000; // 004007c4: LW, REG[3]<=RAM[REG[3]+0];
      10'h1f2: data = 32'h00000000; // 004007c8: SLL, REG[0]<=REG[0]<<0;
      10'h1f3: data = 32'hac430000; // 004007cc: SW, RAM[REG[2]+0]<=REG[3];
      10'h1f4: data = 32'h0810022f; // 004007d0: J, PC<=0x0010022f*4(=0x004008bc);
      10'h1f5: data = 32'h00000000; // 004007d4: SLL, REG[0]<=REG[0]<<0;
      10'h1f6: data = 32'h8fc20008; // 004007d8: LW, REG[2]<=RAM[REG[30]+8];
      10'h1f7: data = 32'h00000000; // 004007dc: SLL, REG[0]<=REG[0]<<0;
      10'h1f8: data = 32'h8c430000; // 004007e0: LW, REG[3]<=RAM[REG[2]+0];
      10'h1f9: data = 32'h2402003f; // 004007e4: ADDIU, REG[2]<=REG[0]+63(=0x0000003f);
      10'h1fa: data = 32'h14620006; // 004007e8: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h1fb: data = 32'h00000000; // 004007ec: SLL, REG[0]<=REG[0]<<0;
      10'h1fc: data = 32'h24030304; // 004007f0: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h1fd: data = 32'h2402003a; // 004007f4: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h1fe: data = 32'hac620000; // 004007f8: SW, RAM[REG[3]+0]<=REG[2];
      10'h1ff: data = 32'h0810022f; // 004007fc: J, PC<=0x0010022f*4(=0x004008bc);
      10'h200: data = 32'h00000000; // 00400800: SLL, REG[0]<=REG[0]<<0;
      10'h201: data = 32'h8fc20008; // 00400804: LW, REG[2]<=RAM[REG[30]+8];
      10'h202: data = 32'h00000000; // 00400808: SLL, REG[0]<=REG[0]<<0;
      10'h203: data = 32'h8c430000; // 0040080c: LW, REG[3]<=RAM[REG[2]+0];
      10'h204: data = 32'h2402003d; // 00400810: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h205: data = 32'h14620006; // 00400814: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h206: data = 32'h00000000; // 00400818: SLL, REG[0]<=REG[0]<<0;
      10'h207: data = 32'h24030304; // 0040081c: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h208: data = 32'h2402003b; // 00400820: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h209: data = 32'hac620000; // 00400824: SW, RAM[REG[3]+0]<=REG[2];
      10'h20a: data = 32'h0810022f; // 00400828: J, PC<=0x0010022f*4(=0x004008bc);
      10'h20b: data = 32'h00000000; // 0040082c: SLL, REG[0]<=REG[0]<<0;
      10'h20c: data = 32'h8fc20008; // 00400830: LW, REG[2]<=RAM[REG[30]+8];
      10'h20d: data = 32'h00000000; // 00400834: SLL, REG[0]<=REG[0]<<0;
      10'h20e: data = 32'h8c430000; // 00400838: LW, REG[3]<=RAM[REG[2]+0];
      10'h20f: data = 32'h2402003b; // 0040083c: ADDIU, REG[2]<=REG[0]+59(=0x0000003b);
      10'h210: data = 32'h14620006; // 00400840: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h211: data = 32'h00000000; // 00400844: SLL, REG[0]<=REG[0]<<0;
      10'h212: data = 32'h24030304; // 00400848: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h213: data = 32'h2402003c; // 0040084c: ADDIU, REG[2]<=REG[0]+60(=0x0000003c);
      10'h214: data = 32'hac620000; // 00400850: SW, RAM[REG[3]+0]<=REG[2];
      10'h215: data = 32'h0810022f; // 00400854: J, PC<=0x0010022f*4(=0x004008bc);
      10'h216: data = 32'h00000000; // 00400858: SLL, REG[0]<=REG[0]<<0;
      10'h217: data = 32'h8fc20008; // 0040085c: LW, REG[2]<=RAM[REG[30]+8];
      10'h218: data = 32'h00000000; // 00400860: SLL, REG[0]<=REG[0]<<0;
      10'h219: data = 32'h8c430000; // 00400864: LW, REG[3]<=RAM[REG[2]+0];
      10'h21a: data = 32'h2402003a; // 00400868: ADDIU, REG[2]<=REG[0]+58(=0x0000003a);
      10'h21b: data = 32'h14620006; // 0040086c: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h21c: data = 32'h00000000; // 00400870: SLL, REG[0]<=REG[0]<<0;
      10'h21d: data = 32'h24030304; // 00400874: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h21e: data = 32'h2402003d; // 00400878: ADDIU, REG[2]<=REG[0]+61(=0x0000003d);
      10'h21f: data = 32'hac620000; // 0040087c: SW, RAM[REG[3]+0]<=REG[2];
      10'h220: data = 32'h0810022f; // 00400880: J, PC<=0x0010022f*4(=0x004008bc);
      10'h221: data = 32'h00000000; // 00400884: SLL, REG[0]<=REG[0]<<0;
      10'h222: data = 32'h8fc20008; // 00400888: LW, REG[2]<=RAM[REG[30]+8];
      10'h223: data = 32'h00000000; // 0040088c: SLL, REG[0]<=REG[0]<<0;
      10'h224: data = 32'h8c430000; // 00400890: LW, REG[3]<=RAM[REG[2]+0];
      10'h225: data = 32'h2402000a; // 00400894: ADDIU, REG[2]<=REG[0]+10(=0x0000000a);
      10'h226: data = 32'h14620006; // 00400898: BNE, PC<=(REG[3] != REG[2])?PC+4+6*4:PC+4;
      10'h227: data = 32'h00000000; // 0040089c: SLL, REG[0]<=REG[0]<<0;
      10'h228: data = 32'h24030304; // 004008a0: ADDIU, REG[3]<=REG[0]+772(=0x00000304);
      10'h229: data = 32'h2402003e; // 004008a4: ADDIU, REG[2]<=REG[0]+62(=0x0000003e);
      10'h22a: data = 32'hac620000; // 004008a8: SW, RAM[REG[3]+0]<=REG[2];
      10'h22b: data = 32'h0810022f; // 004008ac: J, PC<=0x0010022f*4(=0x004008bc);
      10'h22c: data = 32'h00000000; // 004008b0: SLL, REG[0]<=REG[0]<<0;
      10'h22d: data = 32'h24020304; // 004008b4: ADDIU, REG[2]<=REG[0]+772(=0x00000304);
      10'h22e: data = 32'hac400000; // 004008b8: SW, RAM[REG[2]+0]<=REG[0];
      10'h22f: data = 32'h24030300; // 004008bc: ADDIU, REG[3]<=REG[0]+768(=0x00000300);
      10'h230: data = 32'h24020001; // 004008c0: ADDIU, REG[2]<=REG[0]+1(=0x00000001);
      10'h231: data = 32'hac620000; // 004008c4: SW, RAM[REG[3]+0]<=REG[2];
      10'h232: data = 32'h8fc20008; // 004008c8: LW, REG[2]<=RAM[REG[30]+8];
      10'h233: data = 32'h00000000; // 004008cc: SLL, REG[0]<=REG[0]<<0;
      10'h234: data = 32'h24420004; // 004008d0: ADDIU, REG[2]<=REG[2]+4(=0x00000004);
      10'h235: data = 32'hafc20008; // 004008d4: SW, RAM[REG[30]+8]<=REG[2];
      10'h236: data = 32'h8fc20008; // 004008d8: LW, REG[2]<=RAM[REG[30]+8];
      10'h237: data = 32'h00000000; // 004008dc: SLL, REG[0]<=REG[0]<<0;
      10'h238: data = 32'h8c420000; // 004008e0: LW, REG[2]<=RAM[REG[2]+0];
      10'h239: data = 32'h00000000; // 004008e4: SLL, REG[0]<=REG[0]<<0;
      10'h23a: data = 32'h1440ff3f; // 004008e8: BNE, PC<=(REG[2] != REG[0])?PC+4+65343*4:PC+4;
      10'h23b: data = 32'h00000000; // 004008ec: SLL, REG[0]<=REG[0]<<0;
      10'h23c: data = 32'h03c0e821; // 004008f0: ADDU, REG[29]<=REG[30]+REG[0];
      10'h23d: data = 32'h8fbe0000; // 004008f4: LW, REG[30]<=RAM[REG[29]+0];
      10'h23e: data = 32'h27bd0008; // 004008f8: ADDIU, REG[29]<=REG[29]+8(=0x00000008);
      10'h23f: data = 32'h03e00008; // 004008fc: JR, PC<=REG[31];
      10'h240: data = 32'h00000000; // 00400900: SLL, REG[0]<=REG[0]<<0;
      10'h241: data = 32'h27bdfff0; // 00400904: ADDIU, REG[29]<=REG[29]+65520(=0x0000fff0);
      10'h242: data = 32'hafbe0008; // 00400908: SW, RAM[REG[29]+8]<=REG[30];
      10'h243: data = 32'h03a0f021; // 0040090c: ADDU, REG[30]<=REG[29]+REG[0];
      10'h244: data = 32'hafc40010; // 00400910: SW, RAM[REG[30]+16]<=REG[4];
      10'h245: data = 32'h24030320; // 00400914: ADDIU, REG[3]<=REG[0]+800(=0x00000320);
      10'h246: data = 32'h8fc20010; // 00400918: LW, REG[2]<=RAM[REG[30]+16];
      10'h247: data = 32'h00000000; // 0040091c: SLL, REG[0]<=REG[0]<<0;
      10'h248: data = 32'hac620000; // 00400920: SW, RAM[REG[3]+0]<=REG[2];
      10'h249: data = 32'h03c0e821; // 00400924: ADDU, REG[29]<=REG[30]+REG[0];
      10'h24a: data = 32'h8fbe0008; // 00400928: LW, REG[30]<=RAM[REG[29]+8];
      10'h24b: data = 32'h27bd0010; // 0040092c: ADDIU, REG[29]<=REG[29]+16(=0x00000010);
      10'h24c: data = 32'h03e00008; // 00400930: JR, PC<=REG[31];
      10'h24d: data = 32'h00000000; // 00400934: SLL, REG[0]<=REG[0]<<0;
      10'h24e: data = 32'h00000000; // 00400938: SLL, REG[0]<=REG[0]<<0;
      10'h24f: data = 32'h00000000; // 0040093c: SLL, REG[0]<=REG[0]<<0;
    endcase
  end

  assign rom_data = data;
endmodule
